`timescale 1 ns / 1 ns

//yws
module draw_new(clk_25, pause, clk_16, clk_32,clk_8, switchOne, switchTwo, v_count, h_count, rgb, rst, jump);
input               clk_25, clk_16, clk_32,clk_8;
input     [9:0]     v_count;
input     [9:0]     h_count;
input               rst;
input               pause;
input switchOne;
input switchTwo;
input               jump;
output    [7:0]     rgb;
reg       [7:0]     rgb;
   
reg       [9:0]     box_x = 10'd400;
reg       [9:0]     box_y = 10'd200;
parameter [6:0]     box_height = 7'b1001000;
parameter [6:0]     box_width = 7'b1001000;
   
parameter [9:0]     porchleft = 10'b0010010000;   //144
parameter [9:0]     porchtop = 10'b0000100100;    //36
parameter [9:0]     porchbottom = 10'b0111110100; //500
parameter [9:0]     porchright = 10'b1100010000;  //784

parameter BLACK = 8'b000_000_00;
parameter DEFAULT_X = 10'd400;
parameter DEFAULT_Y = 10'd200;
  
reg                 flag_up;
reg                 flag_left;
reg       [5:0]     velocity = 6'd31;   ////pixels/cycle
parameter [5:0] 		velocity_offset  = 6'd31;
                                
reg       [7:0]     accel = 8'd1; //(downwards)
  //6 bits: 0-63

wire [7:0]  rom_dout; 
wire [15:0] addr;
//synthesis attribute box_type <akalin> "black_box" 
//akalin akalin(
//	.clka(clk_25),
//	.addra(addr),
//	.douta(rom_dout)
//	);
assign addr = ((v_count-box_y)*16'd72+(h_count-box_x)); 

reg [31:0] index;
reg frameClk;
reg paused;
initial begin
  paused=0;
  index=0;
end

always @ (*) begin
    if (switchOne) begin
        frameClk = clk_32;
    end
    if (switchTwo) begin
        frameClk = clk_8;
    end
    else begin
        frameClk = clk_16;
    end
end


always @(posedge pause) begin
  paused <= ~paused;
end

always @(posedge frameClk)begin
    //increment index
	 if (paused)begin
		index=index;
	 end
    else if (index==20)begin
      index = 0;
    end
    else
      index = index + 1'b1;
end


always @(posedge clk_25)
begin //DISPLAY
	if(v_count>=36 && v_count<500 && h_count>=144 && h_count<=784)begin
	rgb = frames[index][(v_count-36)/16][(h_count-144)/16];
	end
	else
		rgb=0;
end
   
reg [7:0] frames [0:19][0:29][0:39];	
initial begin
frames[0][0][0] = 8'hb1;
frames[0][0][1] = 8'hb1;
frames[0][0][2] = 8'hb1;
frames[0][0][3] = 8'hd1;
frames[0][0][4] = 8'hd1;
frames[0][0][5] = 8'hd1;
frames[0][0][6] = 8'hd1;
frames[0][0][7] = 8'hd5;
frames[0][0][8] = 8'hd5;
frames[0][0][9] = 8'hd1;
frames[0][0][10] = 8'hd1;
frames[0][0][11] = 8'hd5;
frames[0][0][12] = 8'hd5;
frames[0][0][13] = 8'hd5;
frames[0][0][14] = 8'hd5;
frames[0][0][15] = 8'hd5;
frames[0][0][16] = 8'hd5;
frames[0][0][17] = 8'hd1;
frames[0][0][18] = 8'hd1;
frames[0][0][19] = 8'hd1;
frames[0][0][20] = 8'hd1;
frames[0][0][21] = 8'hd1;
frames[0][0][22] = 8'hd5;
frames[0][0][23] = 8'hd5;
frames[0][0][24] = 8'hd5;
frames[0][0][25] = 8'hd5;
frames[0][0][26] = 8'hd5;
frames[0][0][27] = 8'hd1;
frames[0][0][28] = 8'hd1;
frames[0][0][29] = 8'hd1;
frames[0][0][30] = 8'hd1;
frames[0][0][31] = 8'hd1;
frames[0][0][32] = 8'hd1;
frames[0][0][33] = 8'hd5;
frames[0][0][34] = 8'hd5;
frames[0][0][35] = 8'hd1;
frames[0][0][36] = 8'hd1;
frames[0][0][37] = 8'hd1;
frames[0][0][38] = 8'hb1;
frames[0][0][39] = 8'hb1;
frames[0][1][0] = 8'hb1;
frames[0][1][1] = 8'hb1;
frames[0][1][2] = 8'hb1;
frames[0][1][3] = 8'hd1;
frames[0][1][4] = 8'hd1;
frames[0][1][5] = 8'hd1;
frames[0][1][6] = 8'hd1;
frames[0][1][7] = 8'hd5;
frames[0][1][8] = 8'hd1;
frames[0][1][9] = 8'hd1;
frames[0][1][10] = 8'hd1;
frames[0][1][11] = 8'hd5;
frames[0][1][12] = 8'hd5;
frames[0][1][13] = 8'hd5;
frames[0][1][14] = 8'hd5;
frames[0][1][15] = 8'hd5;
frames[0][1][16] = 8'hd5;
frames[0][1][17] = 8'hd1;
frames[0][1][18] = 8'hd1;
frames[0][1][19] = 8'hd1;
frames[0][1][20] = 8'hd1;
frames[0][1][21] = 8'hd1;
frames[0][1][22] = 8'hd5;
frames[0][1][23] = 8'hd5;
frames[0][1][24] = 8'hd5;
frames[0][1][25] = 8'hd5;
frames[0][1][26] = 8'hd5;
frames[0][1][27] = 8'hd1;
frames[0][1][28] = 8'hd1;
frames[0][1][29] = 8'hd1;
frames[0][1][30] = 8'hd1;
frames[0][1][31] = 8'hd1;
frames[0][1][32] = 8'hd1;
frames[0][1][33] = 8'hd5;
frames[0][1][34] = 8'hd5;
frames[0][1][35] = 8'hd1;
frames[0][1][36] = 8'hd1;
frames[0][1][37] = 8'hd1;
frames[0][1][38] = 8'hb1;
frames[0][1][39] = 8'hb1;
frames[0][2][0] = 8'hb1;
frames[0][2][1] = 8'hb1;
frames[0][2][2] = 8'hd1;
frames[0][2][3] = 8'hd1;
frames[0][2][4] = 8'hd1;
frames[0][2][5] = 8'hd1;
frames[0][2][6] = 8'hd1;
frames[0][2][7] = 8'hd5;
frames[0][2][8] = 8'hd1;
frames[0][2][9] = 8'hd1;
frames[0][2][10] = 8'hd1;
frames[0][2][11] = 8'hd5;
frames[0][2][12] = 8'hd5;
frames[0][2][13] = 8'hd5;
frames[0][2][14] = 8'hd5;
frames[0][2][15] = 8'hd5;
frames[0][2][16] = 8'hd5;
frames[0][2][17] = 8'hd1;
frames[0][2][18] = 8'hd1;
frames[0][2][19] = 8'hd1;
frames[0][2][20] = 8'hd1;
frames[0][2][21] = 8'hd1;
frames[0][2][22] = 8'hd5;
frames[0][2][23] = 8'hd5;
frames[0][2][24] = 8'hd5;
frames[0][2][25] = 8'hd5;
frames[0][2][26] = 8'hd5;
frames[0][2][27] = 8'hd1;
frames[0][2][28] = 8'hd1;
frames[0][2][29] = 8'hd1;
frames[0][2][30] = 8'hd1;
frames[0][2][31] = 8'hd1;
frames[0][2][32] = 8'hd1;
frames[0][2][33] = 8'hd5;
frames[0][2][34] = 8'hd1;
frames[0][2][35] = 8'hd1;
frames[0][2][36] = 8'hd1;
frames[0][2][37] = 8'hd1;
frames[0][2][38] = 8'hb1;
frames[0][2][39] = 8'had;
frames[0][3][0] = 8'hb1;
frames[0][3][1] = 8'hb1;
frames[0][3][2] = 8'hd1;
frames[0][3][3] = 8'hd1;
frames[0][3][4] = 8'hd1;
frames[0][3][5] = 8'hd1;
frames[0][3][6] = 8'hd1;
frames[0][3][7] = 8'hd1;
frames[0][3][8] = 8'hd1;
frames[0][3][9] = 8'hd1;
frames[0][3][10] = 8'hd1;
frames[0][3][11] = 8'hd5;
frames[0][3][12] = 8'hd5;
frames[0][3][13] = 8'hd5;
frames[0][3][14] = 8'hd5;
frames[0][3][15] = 8'hd5;
frames[0][3][16] = 8'hd5;
frames[0][3][17] = 8'hd1;
frames[0][3][18] = 8'hd1;
frames[0][3][19] = 8'hd1;
frames[0][3][20] = 8'hd1;
frames[0][3][21] = 8'hd1;
frames[0][3][22] = 8'hd5;
frames[0][3][23] = 8'hd5;
frames[0][3][24] = 8'hd5;
frames[0][3][25] = 8'hd5;
frames[0][3][26] = 8'hd5;
frames[0][3][27] = 8'hd1;
frames[0][3][28] = 8'hd1;
frames[0][3][29] = 8'hd1;
frames[0][3][30] = 8'hd1;
frames[0][3][31] = 8'hd1;
frames[0][3][32] = 8'hd1;
frames[0][3][33] = 8'hd5;
frames[0][3][34] = 8'hd1;
frames[0][3][35] = 8'hd1;
frames[0][3][36] = 8'hd1;
frames[0][3][37] = 8'hd1;
frames[0][3][38] = 8'hb1;
frames[0][3][39] = 8'had;
frames[0][4][0] = 8'hb1;
frames[0][4][1] = 8'hb1;
frames[0][4][2] = 8'hd1;
frames[0][4][3] = 8'hd1;
frames[0][4][4] = 8'hd1;
frames[0][4][5] = 8'hd1;
frames[0][4][6] = 8'hd1;
frames[0][4][7] = 8'hd1;
frames[0][4][8] = 8'hd1;
frames[0][4][9] = 8'hd1;
frames[0][4][10] = 8'hd1;
frames[0][4][11] = 8'hd5;
frames[0][4][12] = 8'hd5;
frames[0][4][13] = 8'hd5;
frames[0][4][14] = 8'hd5;
frames[0][4][15] = 8'hd5;
frames[0][4][16] = 8'hd5;
frames[0][4][17] = 8'hd1;
frames[0][4][18] = 8'hd1;
frames[0][4][19] = 8'hd1;
frames[0][4][20] = 8'hd1;
frames[0][4][21] = 8'hd1;
frames[0][4][22] = 8'hd5;
frames[0][4][23] = 8'hd5;
frames[0][4][24] = 8'hd5;
frames[0][4][25] = 8'hd5;
frames[0][4][26] = 8'hd5;
frames[0][4][27] = 8'hd5;
frames[0][4][28] = 8'hd1;
frames[0][4][29] = 8'hd1;
frames[0][4][30] = 8'hd1;
frames[0][4][31] = 8'hd1;
frames[0][4][32] = 8'hd1;
frames[0][4][33] = 8'hd5;
frames[0][4][34] = 8'hd1;
frames[0][4][35] = 8'hd1;
frames[0][4][36] = 8'hd1;
frames[0][4][37] = 8'hd1;
frames[0][4][38] = 8'hb1;
frames[0][4][39] = 8'had;
frames[0][5][0] = 8'hb1;
frames[0][5][1] = 8'hb1;
frames[0][5][2] = 8'hd1;
frames[0][5][3] = 8'hd1;
frames[0][5][4] = 8'hd1;
frames[0][5][5] = 8'hd1;
frames[0][5][6] = 8'hd1;
frames[0][5][7] = 8'hd1;
frames[0][5][8] = 8'hd1;
frames[0][5][9] = 8'hd1;
frames[0][5][10] = 8'hd1;
frames[0][5][11] = 8'hd5;
frames[0][5][12] = 8'hd5;
frames[0][5][13] = 8'hd5;
frames[0][5][14] = 8'hd5;
frames[0][5][15] = 8'hd5;
frames[0][5][16] = 8'hd5;
frames[0][5][17] = 8'hd1;
frames[0][5][18] = 8'hd5;
frames[0][5][19] = 8'hd5;
frames[0][5][20] = 8'hd1;
frames[0][5][21] = 8'hd1;
frames[0][5][22] = 8'hd5;
frames[0][5][23] = 8'hd5;
frames[0][5][24] = 8'hd5;
frames[0][5][25] = 8'hd5;
frames[0][5][26] = 8'hd5;
frames[0][5][27] = 8'hd5;
frames[0][5][28] = 8'hd1;
frames[0][5][29] = 8'hd1;
frames[0][5][30] = 8'hd1;
frames[0][5][31] = 8'hd1;
frames[0][5][32] = 8'hd1;
frames[0][5][33] = 8'hd5;
frames[0][5][34] = 8'hd5;
frames[0][5][35] = 8'hd1;
frames[0][5][36] = 8'hd1;
frames[0][5][37] = 8'hd1;
frames[0][5][38] = 8'hd1;
frames[0][5][39] = 8'had;
frames[0][6][0] = 8'hb1;
frames[0][6][1] = 8'hb1;
frames[0][6][2] = 8'hb1;
frames[0][6][3] = 8'hd1;
frames[0][6][4] = 8'hd1;
frames[0][6][5] = 8'hd1;
frames[0][6][6] = 8'hd1;
frames[0][6][7] = 8'hd1;
frames[0][6][8] = 8'hd1;
frames[0][6][9] = 8'hd1;
frames[0][6][10] = 8'hd1;
frames[0][6][11] = 8'hd5;
frames[0][6][12] = 8'hd5;
frames[0][6][13] = 8'hd5;
frames[0][6][14] = 8'hd5;
frames[0][6][15] = 8'hd5;
frames[0][6][16] = 8'hd5;
frames[0][6][17] = 8'hd1;
frames[0][6][18] = 8'hb1;
frames[0][6][19] = 8'h8d;
frames[0][6][20] = 8'h8d;
frames[0][6][21] = 8'hb1;
frames[0][6][22] = 8'hf5;
frames[0][6][23] = 8'hd5;
frames[0][6][24] = 8'hd5;
frames[0][6][25] = 8'hd5;
frames[0][6][26] = 8'hd5;
frames[0][6][27] = 8'hd5;
frames[0][6][28] = 8'hd1;
frames[0][6][29] = 8'hd1;
frames[0][6][30] = 8'hd1;
frames[0][6][31] = 8'hd1;
frames[0][6][32] = 8'hd1;
frames[0][6][33] = 8'hd5;
frames[0][6][34] = 8'hd5;
frames[0][6][35] = 8'hd1;
frames[0][6][36] = 8'hd1;
frames[0][6][37] = 8'hd1;
frames[0][6][38] = 8'hd1;
frames[0][6][39] = 8'had;
frames[0][7][0] = 8'hb1;
frames[0][7][1] = 8'hb1;
frames[0][7][2] = 8'hb1;
frames[0][7][3] = 8'hd1;
frames[0][7][4] = 8'hd1;
frames[0][7][5] = 8'hd1;
frames[0][7][6] = 8'hd1;
frames[0][7][7] = 8'hd1;
frames[0][7][8] = 8'hd1;
frames[0][7][9] = 8'hd1;
frames[0][7][10] = 8'hd1;
frames[0][7][11] = 8'hd5;
frames[0][7][12] = 8'hd5;
frames[0][7][13] = 8'hd5;
frames[0][7][14] = 8'hd5;
frames[0][7][15] = 8'hd5;
frames[0][7][16] = 8'hd5;
frames[0][7][17] = 8'hd1;
frames[0][7][18] = 8'h2a;
frames[0][7][19] = 8'h05;
frames[0][7][20] = 8'h05;
frames[0][7][21] = 8'h2a;
frames[0][7][22] = 8'hd1;
frames[0][7][23] = 8'hd5;
frames[0][7][24] = 8'hd5;
frames[0][7][25] = 8'hd5;
frames[0][7][26] = 8'hd5;
frames[0][7][27] = 8'hd5;
frames[0][7][28] = 8'hd1;
frames[0][7][29] = 8'hd1;
frames[0][7][30] = 8'hd1;
frames[0][7][31] = 8'hd1;
frames[0][7][32] = 8'hd1;
frames[0][7][33] = 8'hd5;
frames[0][7][34] = 8'hd5;
frames[0][7][35] = 8'hd5;
frames[0][7][36] = 8'hd1;
frames[0][7][37] = 8'hd1;
frames[0][7][38] = 8'hd1;
frames[0][7][39] = 8'had;
frames[0][8][0] = 8'hb1;
frames[0][8][1] = 8'hb1;
frames[0][8][2] = 8'hd1;
frames[0][8][3] = 8'hd1;
frames[0][8][4] = 8'hd1;
frames[0][8][5] = 8'hd1;
frames[0][8][6] = 8'hd1;
frames[0][8][7] = 8'hd1;
frames[0][8][8] = 8'hd1;
frames[0][8][9] = 8'hd1;
frames[0][8][10] = 8'hd1;
frames[0][8][11] = 8'hd5;
frames[0][8][12] = 8'hd5;
frames[0][8][13] = 8'hd1;
frames[0][8][14] = 8'hd5;
frames[0][8][15] = 8'hf5;
frames[0][8][16] = 8'hd6;
frames[0][8][17] = 8'h8d;
frames[0][8][18] = 8'h05;
frames[0][8][19] = 8'h05;
frames[0][8][20] = 8'h05;
frames[0][8][21] = 8'h06;
frames[0][8][22] = 8'h91;
frames[0][8][23] = 8'hd6;
frames[0][8][24] = 8'hd5;
frames[0][8][25] = 8'hd5;
frames[0][8][26] = 8'hd5;
frames[0][8][27] = 8'hd5;
frames[0][8][28] = 8'hd5;
frames[0][8][29] = 8'hd5;
frames[0][8][30] = 8'hd1;
frames[0][8][31] = 8'hd1;
frames[0][8][32] = 8'hd1;
frames[0][8][33] = 8'hd5;
frames[0][8][34] = 8'hd5;
frames[0][8][35] = 8'hd5;
frames[0][8][36] = 8'hd1;
frames[0][8][37] = 8'hd1;
frames[0][8][38] = 8'hd1;
frames[0][8][39] = 8'had;
frames[0][9][0] = 8'hb1;
frames[0][9][1] = 8'hb1;
frames[0][9][2] = 8'hd1;
frames[0][9][3] = 8'hd1;
frames[0][9][4] = 8'hd1;
frames[0][9][5] = 8'hd1;
frames[0][9][6] = 8'hd1;
frames[0][9][7] = 8'hd1;
frames[0][9][8] = 8'hd1;
frames[0][9][9] = 8'hd1;
frames[0][9][10] = 8'hd1;
frames[0][9][11] = 8'hd5;
frames[0][9][12] = 8'hd5;
frames[0][9][13] = 8'hd1;
frames[0][9][14] = 8'hd5;
frames[0][9][15] = 8'hf5;
frames[0][9][16] = 8'hd6;
frames[0][9][17] = 8'h8d;
frames[0][9][18] = 8'h4e;
frames[0][9][19] = 8'h4e;
frames[0][9][20] = 8'h73;
frames[0][9][21] = 8'h73;
frames[0][9][22] = 8'h91;
frames[0][9][23] = 8'hd6;
frames[0][9][24] = 8'hd5;
frames[0][9][25] = 8'hd5;
frames[0][9][26] = 8'hd5;
frames[0][9][27] = 8'hd5;
frames[0][9][28] = 8'hd5;
frames[0][9][29] = 8'hd5;
frames[0][9][30] = 8'hd1;
frames[0][9][31] = 8'hd1;
frames[0][9][32] = 8'hd1;
frames[0][9][33] = 8'hd5;
frames[0][9][34] = 8'hd5;
frames[0][9][35] = 8'hd5;
frames[0][9][36] = 8'hd1;
frames[0][9][37] = 8'hd1;
frames[0][9][38] = 8'hd1;
frames[0][9][39] = 8'hb1;
frames[0][10][0] = 8'hb1;
frames[0][10][1] = 8'hb1;
frames[0][10][2] = 8'hd1;
frames[0][10][3] = 8'hd1;
frames[0][10][4] = 8'hd1;
frames[0][10][5] = 8'hd1;
frames[0][10][6] = 8'hd1;
frames[0][10][7] = 8'hd1;
frames[0][10][8] = 8'hd1;
frames[0][10][9] = 8'hd1;
frames[0][10][10] = 8'hd1;
frames[0][10][11] = 8'hd5;
frames[0][10][12] = 8'hd1;
frames[0][10][13] = 8'hd1;
frames[0][10][14] = 8'hd5;
frames[0][10][15] = 8'hf5;
frames[0][10][16] = 8'hd6;
frames[0][10][17] = 8'hb1;
frames[0][10][18] = 8'h93;
frames[0][10][19] = 8'h97;
frames[0][10][20] = 8'h73;
frames[0][10][21] = 8'h2a;
frames[0][10][22] = 8'h6d;
frames[0][10][23] = 8'hd6;
frames[0][10][24] = 8'hd5;
frames[0][10][25] = 8'hd5;
frames[0][10][26] = 8'hd5;
frames[0][10][27] = 8'hd5;
frames[0][10][28] = 8'hd5;
frames[0][10][29] = 8'hd5;
frames[0][10][30] = 8'hd1;
frames[0][10][31] = 8'hd1;
frames[0][10][32] = 8'hd1;
frames[0][10][33] = 8'hd1;
frames[0][10][34] = 8'hd5;
frames[0][10][35] = 8'hd5;
frames[0][10][36] = 8'hd1;
frames[0][10][37] = 8'hd1;
frames[0][10][38] = 8'hd1;
frames[0][10][39] = 8'hb1;
frames[0][11][0] = 8'hb1;
frames[0][11][1] = 8'hb1;
frames[0][11][2] = 8'hd1;
frames[0][11][3] = 8'hd1;
frames[0][11][4] = 8'hd1;
frames[0][11][5] = 8'hd1;
frames[0][11][6] = 8'hd1;
frames[0][11][7] = 8'hd1;
frames[0][11][8] = 8'hd1;
frames[0][11][9] = 8'hd1;
frames[0][11][10] = 8'hd1;
frames[0][11][11] = 8'hd5;
frames[0][11][12] = 8'hd1;
frames[0][11][13] = 8'hd1;
frames[0][11][14] = 8'hd5;
frames[0][11][15] = 8'hf5;
frames[0][11][16] = 8'hd6;
frames[0][11][17] = 8'h8d;
frames[0][11][18] = 8'h2a;
frames[0][11][19] = 8'h0a;
frames[0][11][20] = 8'h05;
frames[0][11][21] = 8'h05;
frames[0][11][22] = 8'h8d;
frames[0][11][23] = 8'hd6;
frames[0][11][24] = 8'hd5;
frames[0][11][25] = 8'hd5;
frames[0][11][26] = 8'hd5;
frames[0][11][27] = 8'hd5;
frames[0][11][28] = 8'hd5;
frames[0][11][29] = 8'hd5;
frames[0][11][30] = 8'hd1;
frames[0][11][31] = 8'hd1;
frames[0][11][32] = 8'hd1;
frames[0][11][33] = 8'hd1;
frames[0][11][34] = 8'hd5;
frames[0][11][35] = 8'hd5;
frames[0][11][36] = 8'hd1;
frames[0][11][37] = 8'hd1;
frames[0][11][38] = 8'hd1;
frames[0][11][39] = 8'hb1;
frames[0][12][0] = 8'had;
frames[0][12][1] = 8'hb1;
frames[0][12][2] = 8'hd1;
frames[0][12][3] = 8'hd1;
frames[0][12][4] = 8'hd1;
frames[0][12][5] = 8'hd1;
frames[0][12][6] = 8'hd1;
frames[0][12][7] = 8'hd1;
frames[0][12][8] = 8'hd1;
frames[0][12][9] = 8'hd1;
frames[0][12][10] = 8'hd1;
frames[0][12][11] = 8'hd5;
frames[0][12][12] = 8'hd1;
frames[0][12][13] = 8'hd1;
frames[0][12][14] = 8'hd5;
frames[0][12][15] = 8'hd5;
frames[0][12][16] = 8'hd5;
frames[0][12][17] = 8'hd1;
frames[0][12][18] = 8'h2a;
frames[0][12][19] = 8'h05;
frames[0][12][20] = 8'h05;
frames[0][12][21] = 8'h2a;
frames[0][12][22] = 8'hd5;
frames[0][12][23] = 8'hd5;
frames[0][12][24] = 8'hd5;
frames[0][12][25] = 8'hd5;
frames[0][12][26] = 8'hf5;
frames[0][12][27] = 8'hd5;
frames[0][12][28] = 8'hd5;
frames[0][12][29] = 8'hd1;
frames[0][12][30] = 8'hd1;
frames[0][12][31] = 8'hd1;
frames[0][12][32] = 8'hd1;
frames[0][12][33] = 8'hd1;
frames[0][12][34] = 8'hd5;
frames[0][12][35] = 8'hd5;
frames[0][12][36] = 8'hd1;
frames[0][12][37] = 8'hd1;
frames[0][12][38] = 8'hd1;
frames[0][12][39] = 8'hb1;
frames[0][13][0] = 8'had;
frames[0][13][1] = 8'hb1;
frames[0][13][2] = 8'hd1;
frames[0][13][3] = 8'hd1;
frames[0][13][4] = 8'hd1;
frames[0][13][5] = 8'hd1;
frames[0][13][6] = 8'hd1;
frames[0][13][7] = 8'hd1;
frames[0][13][8] = 8'hd1;
frames[0][13][9] = 8'hd1;
frames[0][13][10] = 8'hd1;
frames[0][13][11] = 8'hd5;
frames[0][13][12] = 8'hd1;
frames[0][13][13] = 8'hd1;
frames[0][13][14] = 8'hd5;
frames[0][13][15] = 8'hd5;
frames[0][13][16] = 8'hd5;
frames[0][13][17] = 8'hd5;
frames[0][13][18] = 8'hb2;
frames[0][13][19] = 8'h6d;
frames[0][13][20] = 8'h6d;
frames[0][13][21] = 8'h91;
frames[0][13][22] = 8'hd5;
frames[0][13][23] = 8'hd5;
frames[0][13][24] = 8'hd5;
frames[0][13][25] = 8'hd5;
frames[0][13][26] = 8'hd5;
frames[0][13][27] = 8'hd5;
frames[0][13][28] = 8'hd5;
frames[0][13][29] = 8'hd5;
frames[0][13][30] = 8'hd1;
frames[0][13][31] = 8'hd1;
frames[0][13][32] = 8'hd1;
frames[0][13][33] = 8'hd1;
frames[0][13][34] = 8'hd5;
frames[0][13][35] = 8'hd5;
frames[0][13][36] = 8'hd1;
frames[0][13][37] = 8'hd1;
frames[0][13][38] = 8'hb1;
frames[0][13][39] = 8'hb1;
frames[0][14][0] = 8'had;
frames[0][14][1] = 8'hb1;
frames[0][14][2] = 8'hd1;
frames[0][14][3] = 8'hd1;
frames[0][14][4] = 8'hd1;
frames[0][14][5] = 8'hd1;
frames[0][14][6] = 8'hd1;
frames[0][14][7] = 8'hd1;
frames[0][14][8] = 8'hd1;
frames[0][14][9] = 8'hd1;
frames[0][14][10] = 8'hd1;
frames[0][14][11] = 8'hd1;
frames[0][14][12] = 8'hd5;
frames[0][14][13] = 8'hd5;
frames[0][14][14] = 8'hd5;
frames[0][14][15] = 8'hd5;
frames[0][14][16] = 8'hf5;
frames[0][14][17] = 8'hd5;
frames[0][14][18] = 8'hfa;
frames[0][14][19] = 8'hfa;
frames[0][14][20] = 8'hf5;
frames[0][14][21] = 8'hf5;
frames[0][14][22] = 8'hfa;
frames[0][14][23] = 8'hfa;
frames[0][14][24] = 8'hf5;
frames[0][14][25] = 8'hd5;
frames[0][14][26] = 8'hd5;
frames[0][14][27] = 8'hd5;
frames[0][14][28] = 8'hd5;
frames[0][14][29] = 8'hd5;
frames[0][14][30] = 8'hd1;
frames[0][14][31] = 8'hd1;
frames[0][14][32] = 8'hd1;
frames[0][14][33] = 8'hd1;
frames[0][14][34] = 8'hd1;
frames[0][14][35] = 8'hd5;
frames[0][14][36] = 8'hd1;
frames[0][14][37] = 8'hd1;
frames[0][14][38] = 8'hb1;
frames[0][14][39] = 8'hb1;
frames[0][15][0] = 8'had;
frames[0][15][1] = 8'hb1;
frames[0][15][2] = 8'hd1;
frames[0][15][3] = 8'hd1;
frames[0][15][4] = 8'hd1;
frames[0][15][5] = 8'hd1;
frames[0][15][6] = 8'hd1;
frames[0][15][7] = 8'hd1;
frames[0][15][8] = 8'hd1;
frames[0][15][9] = 8'hd1;
frames[0][15][10] = 8'hd1;
frames[0][15][11] = 8'hd1;
frames[0][15][12] = 8'hd5;
frames[0][15][13] = 8'hd5;
frames[0][15][14] = 8'hd5;
frames[0][15][15] = 8'hd5;
frames[0][15][16] = 8'hf6;
frames[0][15][17] = 8'hf6;
frames[0][15][18] = 8'hfa;
frames[0][15][19] = 8'hfa;
frames[0][15][20] = 8'hf6;
frames[0][15][21] = 8'hfa;
frames[0][15][22] = 8'hfa;
frames[0][15][23] = 8'hfa;
frames[0][15][24] = 8'hd5;
frames[0][15][25] = 8'hd5;
frames[0][15][26] = 8'hd5;
frames[0][15][27] = 8'hd5;
frames[0][15][28] = 8'hd5;
frames[0][15][29] = 8'hd5;
frames[0][15][30] = 8'hd1;
frames[0][15][31] = 8'hd1;
frames[0][15][32] = 8'hd1;
frames[0][15][33] = 8'hd1;
frames[0][15][34] = 8'hd1;
frames[0][15][35] = 8'hd1;
frames[0][15][36] = 8'hd1;
frames[0][15][37] = 8'hd1;
frames[0][15][38] = 8'hb1;
frames[0][15][39] = 8'hb1;
frames[0][16][0] = 8'had;
frames[0][16][1] = 8'hb1;
frames[0][16][2] = 8'hb1;
frames[0][16][3] = 8'hb1;
frames[0][16][4] = 8'hd1;
frames[0][16][5] = 8'hd1;
frames[0][16][6] = 8'hd1;
frames[0][16][7] = 8'hd1;
frames[0][16][8] = 8'hd1;
frames[0][16][9] = 8'hd1;
frames[0][16][10] = 8'hd5;
frames[0][16][11] = 8'hd5;
frames[0][16][12] = 8'hd1;
frames[0][16][13] = 8'hd1;
frames[0][16][14] = 8'hd5;
frames[0][16][15] = 8'hf5;
frames[0][16][16] = 8'hd5;
frames[0][16][17] = 8'hd5;
frames[0][16][18] = 8'hd5;
frames[0][16][19] = 8'hf5;
frames[0][16][20] = 8'hd5;
frames[0][16][21] = 8'hd5;
frames[0][16][22] = 8'hf6;
frames[0][16][23] = 8'hf6;
frames[0][16][24] = 8'hf5;
frames[0][16][25] = 8'hd5;
frames[0][16][26] = 8'hd5;
frames[0][16][27] = 8'hd5;
frames[0][16][28] = 8'hd5;
frames[0][16][29] = 8'hd5;
frames[0][16][30] = 8'hd1;
frames[0][16][31] = 8'hd1;
frames[0][16][32] = 8'hd1;
frames[0][16][33] = 8'hd1;
frames[0][16][34] = 8'hd1;
frames[0][16][35] = 8'hd1;
frames[0][16][36] = 8'hd1;
frames[0][16][37] = 8'hb1;
frames[0][16][38] = 8'hb1;
frames[0][16][39] = 8'hb1;
frames[0][17][0] = 8'had;
frames[0][17][1] = 8'hb1;
frames[0][17][2] = 8'hb1;
frames[0][17][3] = 8'hb1;
frames[0][17][4] = 8'hd1;
frames[0][17][5] = 8'hd1;
frames[0][17][6] = 8'hd1;
frames[0][17][7] = 8'hd1;
frames[0][17][8] = 8'hd1;
frames[0][17][9] = 8'hd1;
frames[0][17][10] = 8'hd5;
frames[0][17][11] = 8'hd5;
frames[0][17][12] = 8'hd1;
frames[0][17][13] = 8'hd1;
frames[0][17][14] = 8'hd6;
frames[0][17][15] = 8'hfa;
frames[0][17][16] = 8'hfa;
frames[0][17][17] = 8'hd6;
frames[0][17][18] = 8'hf6;
frames[0][17][19] = 8'hfa;
frames[0][17][20] = 8'hd6;
frames[0][17][21] = 8'hf6;
frames[0][17][22] = 8'hfa;
frames[0][17][23] = 8'hfa;
frames[0][17][24] = 8'hfa;
frames[0][17][25] = 8'hd6;
frames[0][17][26] = 8'hd5;
frames[0][17][27] = 8'hd5;
frames[0][17][28] = 8'hd5;
frames[0][17][29] = 8'hd5;
frames[0][17][30] = 8'hd1;
frames[0][17][31] = 8'hd1;
frames[0][17][32] = 8'hd1;
frames[0][17][33] = 8'hd1;
frames[0][17][34] = 8'hd1;
frames[0][17][35] = 8'hd1;
frames[0][17][36] = 8'hd1;
frames[0][17][37] = 8'hb1;
frames[0][17][38] = 8'hb1;
frames[0][17][39] = 8'hb1;
frames[0][18][0] = 8'had;
frames[0][18][1] = 8'hb1;
frames[0][18][2] = 8'hb1;
frames[0][18][3] = 8'hb1;
frames[0][18][4] = 8'hd1;
frames[0][18][5] = 8'hd1;
frames[0][18][6] = 8'hd1;
frames[0][18][7] = 8'hd1;
frames[0][18][8] = 8'hd1;
frames[0][18][9] = 8'hd1;
frames[0][18][10] = 8'hd5;
frames[0][18][11] = 8'hd5;
frames[0][18][12] = 8'hd5;
frames[0][18][13] = 8'hd1;
frames[0][18][14] = 8'hd6;
frames[0][18][15] = 8'hfa;
frames[0][18][16] = 8'hfa;
frames[0][18][17] = 8'hd6;
frames[0][18][18] = 8'hf6;
frames[0][18][19] = 8'hfa;
frames[0][18][20] = 8'hd6;
frames[0][18][21] = 8'hfa;
frames[0][18][22] = 8'hfa;
frames[0][18][23] = 8'hd6;
frames[0][18][24] = 8'hfa;
frames[0][18][25] = 8'hf6;
frames[0][18][26] = 8'hd5;
frames[0][18][27] = 8'hd5;
frames[0][18][28] = 8'hd5;
frames[0][18][29] = 8'hd1;
frames[0][18][30] = 8'hd1;
frames[0][18][31] = 8'hd1;
frames[0][18][32] = 8'hd1;
frames[0][18][33] = 8'hd1;
frames[0][18][34] = 8'hd1;
frames[0][18][35] = 8'hd1;
frames[0][18][36] = 8'hd1;
frames[0][18][37] = 8'hb1;
frames[0][18][38] = 8'hb1;
frames[0][18][39] = 8'hb1;
frames[0][19][0] = 8'hac;
frames[0][19][1] = 8'hb1;
frames[0][19][2] = 8'hb1;
frames[0][19][3] = 8'hb1;
frames[0][19][4] = 8'hd1;
frames[0][19][5] = 8'hd1;
frames[0][19][6] = 8'hd1;
frames[0][19][7] = 8'hd1;
frames[0][19][8] = 8'hd1;
frames[0][19][9] = 8'hd1;
frames[0][19][10] = 8'hd5;
frames[0][19][11] = 8'hd5;
frames[0][19][12] = 8'hd5;
frames[0][19][13] = 8'hd1;
frames[0][19][14] = 8'hd6;
frames[0][19][15] = 8'hfa;
frames[0][19][16] = 8'hfa;
frames[0][19][17] = 8'hda;
frames[0][19][18] = 8'hfa;
frames[0][19][19] = 8'hfa;
frames[0][19][20] = 8'hd5;
frames[0][19][21] = 8'hd5;
frames[0][19][22] = 8'hfa;
frames[0][19][23] = 8'hfa;
frames[0][19][24] = 8'hfa;
frames[0][19][25] = 8'hd6;
frames[0][19][26] = 8'hd5;
frames[0][19][27] = 8'hd5;
frames[0][19][28] = 8'hd1;
frames[0][19][29] = 8'hd1;
frames[0][19][30] = 8'hd1;
frames[0][19][31] = 8'hd1;
frames[0][19][32] = 8'hd1;
frames[0][19][33] = 8'hd1;
frames[0][19][34] = 8'hd1;
frames[0][19][35] = 8'hd1;
frames[0][19][36] = 8'hd1;
frames[0][19][37] = 8'hb1;
frames[0][19][38] = 8'hb1;
frames[0][19][39] = 8'hb1;
frames[0][20][0] = 8'hac;
frames[0][20][1] = 8'hb1;
frames[0][20][2] = 8'hb1;
frames[0][20][3] = 8'hb1;
frames[0][20][4] = 8'hd1;
frames[0][20][5] = 8'hd1;
frames[0][20][6] = 8'hd1;
frames[0][20][7] = 8'hd1;
frames[0][20][8] = 8'hd1;
frames[0][20][9] = 8'hd1;
frames[0][20][10] = 8'hd5;
frames[0][20][11] = 8'hd5;
frames[0][20][12] = 8'hd5;
frames[0][20][13] = 8'hd5;
frames[0][20][14] = 8'hd5;
frames[0][20][15] = 8'hf5;
frames[0][20][16] = 8'hd5;
frames[0][20][17] = 8'hf6;
frames[0][20][18] = 8'hf6;
frames[0][20][19] = 8'hf6;
frames[0][20][20] = 8'hd5;
frames[0][20][21] = 8'hd5;
frames[0][20][22] = 8'hd6;
frames[0][20][23] = 8'hf6;
frames[0][20][24] = 8'hf6;
frames[0][20][25] = 8'hd5;
frames[0][20][26] = 8'hd5;
frames[0][20][27] = 8'hd5;
frames[0][20][28] = 8'hd5;
frames[0][20][29] = 8'hd1;
frames[0][20][30] = 8'hd1;
frames[0][20][31] = 8'hd1;
frames[0][20][32] = 8'hd1;
frames[0][20][33] = 8'hd1;
frames[0][20][34] = 8'hd1;
frames[0][20][35] = 8'hd1;
frames[0][20][36] = 8'hb1;
frames[0][20][37] = 8'hb1;
frames[0][20][38] = 8'hb1;
frames[0][20][39] = 8'hb1;
frames[0][21][0] = 8'hac;
frames[0][21][1] = 8'hb1;
frames[0][21][2] = 8'hb1;
frames[0][21][3] = 8'hb1;
frames[0][21][4] = 8'hd1;
frames[0][21][5] = 8'hd1;
frames[0][21][6] = 8'hd1;
frames[0][21][7] = 8'hd1;
frames[0][21][8] = 8'hd1;
frames[0][21][9] = 8'hd1;
frames[0][21][10] = 8'hd1;
frames[0][21][11] = 8'hd1;
frames[0][21][12] = 8'hd5;
frames[0][21][13] = 8'hd5;
frames[0][21][14] = 8'hd5;
frames[0][21][15] = 8'hf6;
frames[0][21][16] = 8'hfa;
frames[0][21][17] = 8'hfa;
frames[0][21][18] = 8'hfa;
frames[0][21][19] = 8'hfa;
frames[0][21][20] = 8'hfa;
frames[0][21][21] = 8'hf6;
frames[0][21][22] = 8'hd6;
frames[0][21][23] = 8'hfa;
frames[0][21][24] = 8'hf6;
frames[0][21][25] = 8'hd5;
frames[0][21][26] = 8'hd5;
frames[0][21][27] = 8'hd5;
frames[0][21][28] = 8'hd5;
frames[0][21][29] = 8'hd1;
frames[0][21][30] = 8'hd1;
frames[0][21][31] = 8'hd1;
frames[0][21][32] = 8'hd1;
frames[0][21][33] = 8'hd1;
frames[0][21][34] = 8'hb1;
frames[0][21][35] = 8'hd1;
frames[0][21][36] = 8'hb1;
frames[0][21][37] = 8'hb1;
frames[0][21][38] = 8'hb1;
frames[0][21][39] = 8'hb1;
frames[0][22][0] = 8'hac;
frames[0][22][1] = 8'hb1;
frames[0][22][2] = 8'hb1;
frames[0][22][3] = 8'hb1;
frames[0][22][4] = 8'hb1;
frames[0][22][5] = 8'hd1;
frames[0][22][6] = 8'hd1;
frames[0][22][7] = 8'hd1;
frames[0][22][8] = 8'hd1;
frames[0][22][9] = 8'hd1;
frames[0][22][10] = 8'hd1;
frames[0][22][11] = 8'hd1;
frames[0][22][12] = 8'hd5;
frames[0][22][13] = 8'hd5;
frames[0][22][14] = 8'hd5;
frames[0][22][15] = 8'hf6;
frames[0][22][16] = 8'hfa;
frames[0][22][17] = 8'hfa;
frames[0][22][18] = 8'hd6;
frames[0][22][19] = 8'hfa;
frames[0][22][20] = 8'hfa;
frames[0][22][21] = 8'hfa;
frames[0][22][22] = 8'hd6;
frames[0][22][23] = 8'hfa;
frames[0][22][24] = 8'hf6;
frames[0][22][25] = 8'hd5;
frames[0][22][26] = 8'hd5;
frames[0][22][27] = 8'hd1;
frames[0][22][28] = 8'hd1;
frames[0][22][29] = 8'hd1;
frames[0][22][30] = 8'hd1;
frames[0][22][31] = 8'hd1;
frames[0][22][32] = 8'hd1;
frames[0][22][33] = 8'hd1;
frames[0][22][34] = 8'hb1;
frames[0][22][35] = 8'hd1;
frames[0][22][36] = 8'hb1;
frames[0][22][37] = 8'hb1;
frames[0][22][38] = 8'hb1;
frames[0][22][39] = 8'hb1;
frames[0][23][0] = 8'hac;
frames[0][23][1] = 8'hb1;
frames[0][23][2] = 8'hb1;
frames[0][23][3] = 8'hb1;
frames[0][23][4] = 8'hb1;
frames[0][23][5] = 8'hd1;
frames[0][23][6] = 8'hd1;
frames[0][23][7] = 8'hd1;
frames[0][23][8] = 8'hd1;
frames[0][23][9] = 8'hd1;
frames[0][23][10] = 8'hd1;
frames[0][23][11] = 8'hd1;
frames[0][23][12] = 8'hd1;
frames[0][23][13] = 8'hd5;
frames[0][23][14] = 8'hd5;
frames[0][23][15] = 8'hfa;
frames[0][23][16] = 8'hfa;
frames[0][23][17] = 8'hfa;
frames[0][23][18] = 8'hfa;
frames[0][23][19] = 8'hfa;
frames[0][23][20] = 8'hfa;
frames[0][23][21] = 8'hfa;
frames[0][23][22] = 8'hfa;
frames[0][23][23] = 8'hfa;
frames[0][23][24] = 8'hfa;
frames[0][23][25] = 8'hd5;
frames[0][23][26] = 8'hd1;
frames[0][23][27] = 8'hd1;
frames[0][23][28] = 8'hd1;
frames[0][23][29] = 8'hd1;
frames[0][23][30] = 8'hd1;
frames[0][23][31] = 8'hd1;
frames[0][23][32] = 8'hd1;
frames[0][23][33] = 8'hb1;
frames[0][23][34] = 8'hb1;
frames[0][23][35] = 8'hd1;
frames[0][23][36] = 8'hb1;
frames[0][23][37] = 8'hb1;
frames[0][23][38] = 8'hb1;
frames[0][23][39] = 8'hb1;
frames[0][24][0] = 8'hac;
frames[0][24][1] = 8'hb1;
frames[0][24][2] = 8'hb1;
frames[0][24][3] = 8'hb1;
frames[0][24][4] = 8'hb1;
frames[0][24][5] = 8'hd1;
frames[0][24][6] = 8'hd1;
frames[0][24][7] = 8'hd1;
frames[0][24][8] = 8'hd1;
frames[0][24][9] = 8'hd1;
frames[0][24][10] = 8'hd1;
frames[0][24][11] = 8'hd1;
frames[0][24][12] = 8'hd1;
frames[0][24][13] = 8'hd1;
frames[0][24][14] = 8'hd5;
frames[0][24][15] = 8'hd5;
frames[0][24][16] = 8'hd5;
frames[0][24][17] = 8'hd5;
frames[0][24][18] = 8'hd5;
frames[0][24][19] = 8'hd5;
frames[0][24][20] = 8'hd5;
frames[0][24][21] = 8'hd5;
frames[0][24][22] = 8'hd5;
frames[0][24][23] = 8'hd5;
frames[0][24][24] = 8'hd5;
frames[0][24][25] = 8'hd5;
frames[0][24][26] = 8'hd1;
frames[0][24][27] = 8'hd1;
frames[0][24][28] = 8'hd1;
frames[0][24][29] = 8'hd1;
frames[0][24][30] = 8'hd1;
frames[0][24][31] = 8'hd1;
frames[0][24][32] = 8'hb1;
frames[0][24][33] = 8'hb1;
frames[0][24][34] = 8'hb1;
frames[0][24][35] = 8'hd1;
frames[0][24][36] = 8'hb1;
frames[0][24][37] = 8'hb1;
frames[0][24][38] = 8'hb1;
frames[0][24][39] = 8'hb1;
frames[0][25][0] = 8'hac;
frames[0][25][1] = 8'hac;
frames[0][25][2] = 8'hac;
frames[0][25][3] = 8'hac;
frames[0][25][4] = 8'hb1;
frames[0][25][5] = 8'hd1;
frames[0][25][6] = 8'hd1;
frames[0][25][7] = 8'hd1;
frames[0][25][8] = 8'hd1;
frames[0][25][9] = 8'hd1;
frames[0][25][10] = 8'hd1;
frames[0][25][11] = 8'hd1;
frames[0][25][12] = 8'hd1;
frames[0][25][13] = 8'hd1;
frames[0][25][14] = 8'hd1;
frames[0][25][15] = 8'hd1;
frames[0][25][16] = 8'hd1;
frames[0][25][17] = 8'hd1;
frames[0][25][18] = 8'hd1;
frames[0][25][19] = 8'hd5;
frames[0][25][20] = 8'hd5;
frames[0][25][21] = 8'hd5;
frames[0][25][22] = 8'hd5;
frames[0][25][23] = 8'hd5;
frames[0][25][24] = 8'hd5;
frames[0][25][25] = 8'hd5;
frames[0][25][26] = 8'hd1;
frames[0][25][27] = 8'hd1;
frames[0][25][28] = 8'hd1;
frames[0][25][29] = 8'hd1;
frames[0][25][30] = 8'hd1;
frames[0][25][31] = 8'hd1;
frames[0][25][32] = 8'hb1;
frames[0][25][33] = 8'hb1;
frames[0][25][34] = 8'hb1;
frames[0][25][35] = 8'hb1;
frames[0][25][36] = 8'hb1;
frames[0][25][37] = 8'hb1;
frames[0][25][38] = 8'hb1;
frames[0][25][39] = 8'hb1;
frames[0][26][0] = 8'h8c;
frames[0][26][1] = 8'hac;
frames[0][26][2] = 8'hac;
frames[0][26][3] = 8'hac;
frames[0][26][4] = 8'hb0;
frames[0][26][5] = 8'hb1;
frames[0][26][6] = 8'hd1;
frames[0][26][7] = 8'hd1;
frames[0][26][8] = 8'hd1;
frames[0][26][9] = 8'hd1;
frames[0][26][10] = 8'hd1;
frames[0][26][11] = 8'hd1;
frames[0][26][12] = 8'hd1;
frames[0][26][13] = 8'hd1;
frames[0][26][14] = 8'hd1;
frames[0][26][15] = 8'hd1;
frames[0][26][16] = 8'hd1;
frames[0][26][17] = 8'hd1;
frames[0][26][18] = 8'hd1;
frames[0][26][19] = 8'hd1;
frames[0][26][20] = 8'hd1;
frames[0][26][21] = 8'hd1;
frames[0][26][22] = 8'hd5;
frames[0][26][23] = 8'hd5;
frames[0][26][24] = 8'hd5;
frames[0][26][25] = 8'hd1;
frames[0][26][26] = 8'hd1;
frames[0][26][27] = 8'hd1;
frames[0][26][28] = 8'hd1;
frames[0][26][29] = 8'hd1;
frames[0][26][30] = 8'hd1;
frames[0][26][31] = 8'hb1;
frames[0][26][32] = 8'hb1;
frames[0][26][33] = 8'hb1;
frames[0][26][34] = 8'hb1;
frames[0][26][35] = 8'hb1;
frames[0][26][36] = 8'hb1;
frames[0][26][37] = 8'hb1;
frames[0][26][38] = 8'hb1;
frames[0][26][39] = 8'hb1;
frames[0][27][0] = 8'h8c;
frames[0][27][1] = 8'hac;
frames[0][27][2] = 8'hac;
frames[0][27][3] = 8'hac;
frames[0][27][4] = 8'hac;
frames[0][27][5] = 8'hb1;
frames[0][27][6] = 8'hd1;
frames[0][27][7] = 8'hd1;
frames[0][27][8] = 8'hd1;
frames[0][27][9] = 8'hd1;
frames[0][27][10] = 8'hd1;
frames[0][27][11] = 8'hd1;
frames[0][27][12] = 8'hd1;
frames[0][27][13] = 8'hd1;
frames[0][27][14] = 8'hd1;
frames[0][27][15] = 8'hd1;
frames[0][27][16] = 8'hb1;
frames[0][27][17] = 8'hb1;
frames[0][27][18] = 8'hb1;
frames[0][27][19] = 8'hd1;
frames[0][27][20] = 8'hd1;
frames[0][27][21] = 8'hd1;
frames[0][27][22] = 8'hd1;
frames[0][27][23] = 8'hd1;
frames[0][27][24] = 8'hd1;
frames[0][27][25] = 8'hd1;
frames[0][27][26] = 8'hd1;
frames[0][27][27] = 8'hd1;
frames[0][27][28] = 8'hd1;
frames[0][27][29] = 8'hd1;
frames[0][27][30] = 8'hd1;
frames[0][27][31] = 8'hb1;
frames[0][27][32] = 8'hb1;
frames[0][27][33] = 8'hb1;
frames[0][27][34] = 8'hb1;
frames[0][27][35] = 8'hb1;
frames[0][27][36] = 8'hb1;
frames[0][27][37] = 8'hb1;
frames[0][27][38] = 8'hb1;
frames[0][27][39] = 8'hb1;
frames[0][28][0] = 8'h8c;
frames[0][28][1] = 8'h8c;
frames[0][28][2] = 8'h8c;
frames[0][28][3] = 8'hac;
frames[0][28][4] = 8'hac;
frames[0][28][5] = 8'had;
frames[0][28][6] = 8'hb1;
frames[0][28][7] = 8'hb1;
frames[0][28][8] = 8'hd1;
frames[0][28][9] = 8'hd1;
frames[0][28][10] = 8'hd1;
frames[0][28][11] = 8'hd1;
frames[0][28][12] = 8'hd1;
frames[0][28][13] = 8'hd1;
frames[0][28][14] = 8'hd1;
frames[0][28][15] = 8'hd1;
frames[0][28][16] = 8'had;
frames[0][28][17] = 8'hac;
frames[0][28][18] = 8'had;
frames[0][28][19] = 8'had;
frames[0][28][20] = 8'hb1;
frames[0][28][21] = 8'hb1;
frames[0][28][22] = 8'hd1;
frames[0][28][23] = 8'hd1;
frames[0][28][24] = 8'hd1;
frames[0][28][25] = 8'hd1;
frames[0][28][26] = 8'hd1;
frames[0][28][27] = 8'hb1;
frames[0][28][28] = 8'hb1;
frames[0][28][29] = 8'hb1;
frames[0][28][30] = 8'hb1;
frames[0][28][31] = 8'hb1;
frames[0][28][32] = 8'hb1;
frames[0][28][33] = 8'hb1;
frames[0][28][34] = 8'hb1;
frames[0][28][35] = 8'hb1;
frames[0][28][36] = 8'hb1;
frames[0][28][37] = 8'hb1;
frames[0][28][38] = 8'hb1;
frames[0][28][39] = 8'had;
frames[0][29][0] = 8'h8c;
frames[0][29][1] = 8'h8c;
frames[0][29][2] = 8'h8c;
frames[0][29][3] = 8'h8c;
frames[0][29][4] = 8'hac;
frames[0][29][5] = 8'hac;
frames[0][29][6] = 8'hac;
frames[0][29][7] = 8'hb1;
frames[0][29][8] = 8'hd1;
frames[0][29][9] = 8'hd1;
frames[0][29][10] = 8'hd1;
frames[0][29][11] = 8'hd1;
frames[0][29][12] = 8'hd1;
frames[0][29][13] = 8'hd1;
frames[0][29][14] = 8'hd1;
frames[0][29][15] = 8'hd1;
frames[0][29][16] = 8'had;
frames[0][29][17] = 8'hac;
frames[0][29][18] = 8'hac;
frames[0][29][19] = 8'hac;
frames[0][29][20] = 8'hac;
frames[0][29][21] = 8'hac;
frames[0][29][22] = 8'hb1;
frames[0][29][23] = 8'hd1;
frames[0][29][24] = 8'hd1;
frames[0][29][25] = 8'hd1;
frames[0][29][26] = 8'hb1;
frames[0][29][27] = 8'hb1;
frames[0][29][28] = 8'hb1;
frames[0][29][29] = 8'hb1;
frames[0][29][30] = 8'hb1;
frames[0][29][31] = 8'hb1;
frames[0][29][32] = 8'hb1;
frames[0][29][33] = 8'hb1;
frames[0][29][34] = 8'hb1;
frames[0][29][35] = 8'hb1;
frames[0][29][36] = 8'hb1;
frames[0][29][37] = 8'hb1;
frames[0][29][38] = 8'hb1;
frames[0][29][39] = 8'hb1;
frames[1][0][0] = 8'hb1;
frames[1][0][1] = 8'hb1;
frames[1][0][2] = 8'hb1;
frames[1][0][3] = 8'hd1;
frames[1][0][4] = 8'hd1;
frames[1][0][5] = 8'hd1;
frames[1][0][6] = 8'hd1;
frames[1][0][7] = 8'hd5;
frames[1][0][8] = 8'hd5;
frames[1][0][9] = 8'hd1;
frames[1][0][10] = 8'hd1;
frames[1][0][11] = 8'hd5;
frames[1][0][12] = 8'hd5;
frames[1][0][13] = 8'hd5;
frames[1][0][14] = 8'hd5;
frames[1][0][15] = 8'hd5;
frames[1][0][16] = 8'hd5;
frames[1][0][17] = 8'hd1;
frames[1][0][18] = 8'hd1;
frames[1][0][19] = 8'hd1;
frames[1][0][20] = 8'hd1;
frames[1][0][21] = 8'hd1;
frames[1][0][22] = 8'hd5;
frames[1][0][23] = 8'hd5;
frames[1][0][24] = 8'hd5;
frames[1][0][25] = 8'hd5;
frames[1][0][26] = 8'hd5;
frames[1][0][27] = 8'hd1;
frames[1][0][28] = 8'hd1;
frames[1][0][29] = 8'hd1;
frames[1][0][30] = 8'hd1;
frames[1][0][31] = 8'hd1;
frames[1][0][32] = 8'hd1;
frames[1][0][33] = 8'hd5;
frames[1][0][34] = 8'hd5;
frames[1][0][35] = 8'hd1;
frames[1][0][36] = 8'hd1;
frames[1][0][37] = 8'hd1;
frames[1][0][38] = 8'hb1;
frames[1][0][39] = 8'hb1;
frames[1][1][0] = 8'hb1;
frames[1][1][1] = 8'hb1;
frames[1][1][2] = 8'hb1;
frames[1][1][3] = 8'hd1;
frames[1][1][4] = 8'hd1;
frames[1][1][5] = 8'hd1;
frames[1][1][6] = 8'hd1;
frames[1][1][7] = 8'hd5;
frames[1][1][8] = 8'hd1;
frames[1][1][9] = 8'hd1;
frames[1][1][10] = 8'hd1;
frames[1][1][11] = 8'hd5;
frames[1][1][12] = 8'hd5;
frames[1][1][13] = 8'hd5;
frames[1][1][14] = 8'hd5;
frames[1][1][15] = 8'hd5;
frames[1][1][16] = 8'hd5;
frames[1][1][17] = 8'hd1;
frames[1][1][18] = 8'hd1;
frames[1][1][19] = 8'hd1;
frames[1][1][20] = 8'hd1;
frames[1][1][21] = 8'hd1;
frames[1][1][22] = 8'hd5;
frames[1][1][23] = 8'hd5;
frames[1][1][24] = 8'hd5;
frames[1][1][25] = 8'hd5;
frames[1][1][26] = 8'hd5;
frames[1][1][27] = 8'hd1;
frames[1][1][28] = 8'hd1;
frames[1][1][29] = 8'hd1;
frames[1][1][30] = 8'hd1;
frames[1][1][31] = 8'hd1;
frames[1][1][32] = 8'hd1;
frames[1][1][33] = 8'hd5;
frames[1][1][34] = 8'hd5;
frames[1][1][35] = 8'hd1;
frames[1][1][36] = 8'hd1;
frames[1][1][37] = 8'hd1;
frames[1][1][38] = 8'hb1;
frames[1][1][39] = 8'hb1;
frames[1][2][0] = 8'hb1;
frames[1][2][1] = 8'hb1;
frames[1][2][2] = 8'hd1;
frames[1][2][3] = 8'hd1;
frames[1][2][4] = 8'hd1;
frames[1][2][5] = 8'hd1;
frames[1][2][6] = 8'hd1;
frames[1][2][7] = 8'hd5;
frames[1][2][8] = 8'hd1;
frames[1][2][9] = 8'hd1;
frames[1][2][10] = 8'hd1;
frames[1][2][11] = 8'hd5;
frames[1][2][12] = 8'hd5;
frames[1][2][13] = 8'hd5;
frames[1][2][14] = 8'hd5;
frames[1][2][15] = 8'hd5;
frames[1][2][16] = 8'hd5;
frames[1][2][17] = 8'hd1;
frames[1][2][18] = 8'hd1;
frames[1][2][19] = 8'hd1;
frames[1][2][20] = 8'hd1;
frames[1][2][21] = 8'hd1;
frames[1][2][22] = 8'hd5;
frames[1][2][23] = 8'hd5;
frames[1][2][24] = 8'hd5;
frames[1][2][25] = 8'hd5;
frames[1][2][26] = 8'hd5;
frames[1][2][27] = 8'hd1;
frames[1][2][28] = 8'hd1;
frames[1][2][29] = 8'hd1;
frames[1][2][30] = 8'hd1;
frames[1][2][31] = 8'hd1;
frames[1][2][32] = 8'hd1;
frames[1][2][33] = 8'hd5;
frames[1][2][34] = 8'hd1;
frames[1][2][35] = 8'hd1;
frames[1][2][36] = 8'hd1;
frames[1][2][37] = 8'hd1;
frames[1][2][38] = 8'hb1;
frames[1][2][39] = 8'had;
frames[1][3][0] = 8'hb1;
frames[1][3][1] = 8'hb1;
frames[1][3][2] = 8'hd1;
frames[1][3][3] = 8'hd1;
frames[1][3][4] = 8'hd1;
frames[1][3][5] = 8'hd1;
frames[1][3][6] = 8'hd1;
frames[1][3][7] = 8'hd1;
frames[1][3][8] = 8'hd1;
frames[1][3][9] = 8'hd1;
frames[1][3][10] = 8'hd1;
frames[1][3][11] = 8'hd5;
frames[1][3][12] = 8'hd5;
frames[1][3][13] = 8'hd5;
frames[1][3][14] = 8'hd5;
frames[1][3][15] = 8'hd5;
frames[1][3][16] = 8'hd5;
frames[1][3][17] = 8'hd1;
frames[1][3][18] = 8'hd1;
frames[1][3][19] = 8'hd1;
frames[1][3][20] = 8'hd1;
frames[1][3][21] = 8'hd1;
frames[1][3][22] = 8'hd5;
frames[1][3][23] = 8'hd5;
frames[1][3][24] = 8'hd5;
frames[1][3][25] = 8'hd5;
frames[1][3][26] = 8'hd5;
frames[1][3][27] = 8'hd1;
frames[1][3][28] = 8'hd1;
frames[1][3][29] = 8'hd1;
frames[1][3][30] = 8'hd1;
frames[1][3][31] = 8'hd1;
frames[1][3][32] = 8'hd1;
frames[1][3][33] = 8'hd5;
frames[1][3][34] = 8'hd1;
frames[1][3][35] = 8'hd1;
frames[1][3][36] = 8'hd1;
frames[1][3][37] = 8'hd1;
frames[1][3][38] = 8'hb1;
frames[1][3][39] = 8'had;
frames[1][4][0] = 8'hb1;
frames[1][4][1] = 8'hb1;
frames[1][4][2] = 8'hd1;
frames[1][4][3] = 8'hd1;
frames[1][4][4] = 8'hd1;
frames[1][4][5] = 8'hd1;
frames[1][4][6] = 8'hd1;
frames[1][4][7] = 8'hd1;
frames[1][4][8] = 8'hd1;
frames[1][4][9] = 8'hd1;
frames[1][4][10] = 8'hd1;
frames[1][4][11] = 8'hd5;
frames[1][4][12] = 8'hd5;
frames[1][4][13] = 8'hd5;
frames[1][4][14] = 8'hd5;
frames[1][4][15] = 8'hd5;
frames[1][4][16] = 8'hd5;
frames[1][4][17] = 8'hd1;
frames[1][4][18] = 8'hd1;
frames[1][4][19] = 8'hd1;
frames[1][4][20] = 8'hd1;
frames[1][4][21] = 8'hd1;
frames[1][4][22] = 8'hd5;
frames[1][4][23] = 8'hd5;
frames[1][4][24] = 8'hd5;
frames[1][4][25] = 8'hd5;
frames[1][4][26] = 8'hd5;
frames[1][4][27] = 8'hd5;
frames[1][4][28] = 8'hd1;
frames[1][4][29] = 8'hd1;
frames[1][4][30] = 8'hd1;
frames[1][4][31] = 8'hd1;
frames[1][4][32] = 8'hd1;
frames[1][4][33] = 8'hd5;
frames[1][4][34] = 8'hd1;
frames[1][4][35] = 8'hd1;
frames[1][4][36] = 8'hd1;
frames[1][4][37] = 8'hd1;
frames[1][4][38] = 8'hb1;
frames[1][4][39] = 8'had;
frames[1][5][0] = 8'hb1;
frames[1][5][1] = 8'hb1;
frames[1][5][2] = 8'hd1;
frames[1][5][3] = 8'hd1;
frames[1][5][4] = 8'hd1;
frames[1][5][5] = 8'hd1;
frames[1][5][6] = 8'hd1;
frames[1][5][7] = 8'hd1;
frames[1][5][8] = 8'hd1;
frames[1][5][9] = 8'hd1;
frames[1][5][10] = 8'hd1;
frames[1][5][11] = 8'hd5;
frames[1][5][12] = 8'hd5;
frames[1][5][13] = 8'hd5;
frames[1][5][14] = 8'hd5;
frames[1][5][15] = 8'hd5;
frames[1][5][16] = 8'hd5;
frames[1][5][17] = 8'hd1;
frames[1][5][18] = 8'hd5;
frames[1][5][19] = 8'hd5;
frames[1][5][20] = 8'hd1;
frames[1][5][21] = 8'hd1;
frames[1][5][22] = 8'hd5;
frames[1][5][23] = 8'hd5;
frames[1][5][24] = 8'hd5;
frames[1][5][25] = 8'hd5;
frames[1][5][26] = 8'hd5;
frames[1][5][27] = 8'hd5;
frames[1][5][28] = 8'hd1;
frames[1][5][29] = 8'hd1;
frames[1][5][30] = 8'hd1;
frames[1][5][31] = 8'hd1;
frames[1][5][32] = 8'hd1;
frames[1][5][33] = 8'hd5;
frames[1][5][34] = 8'hd5;
frames[1][5][35] = 8'hd1;
frames[1][5][36] = 8'hd1;
frames[1][5][37] = 8'hd1;
frames[1][5][38] = 8'hd1;
frames[1][5][39] = 8'had;
frames[1][6][0] = 8'hb1;
frames[1][6][1] = 8'hb1;
frames[1][6][2] = 8'hb1;
frames[1][6][3] = 8'hd1;
frames[1][6][4] = 8'hd1;
frames[1][6][5] = 8'hd1;
frames[1][6][6] = 8'hd1;
frames[1][6][7] = 8'hd1;
frames[1][6][8] = 8'hd1;
frames[1][6][9] = 8'hd1;
frames[1][6][10] = 8'hd1;
frames[1][6][11] = 8'hd5;
frames[1][6][12] = 8'hd5;
frames[1][6][13] = 8'hd5;
frames[1][6][14] = 8'hd5;
frames[1][6][15] = 8'hd5;
frames[1][6][16] = 8'hd5;
frames[1][6][17] = 8'hd5;
frames[1][6][18] = 8'hb1;
frames[1][6][19] = 8'h8d;
frames[1][6][20] = 8'h8d;
frames[1][6][21] = 8'hb1;
frames[1][6][22] = 8'hf5;
frames[1][6][23] = 8'hd5;
frames[1][6][24] = 8'hd5;
frames[1][6][25] = 8'hd5;
frames[1][6][26] = 8'hd5;
frames[1][6][27] = 8'hd5;
frames[1][6][28] = 8'hd1;
frames[1][6][29] = 8'hd1;
frames[1][6][30] = 8'hd1;
frames[1][6][31] = 8'hd1;
frames[1][6][32] = 8'hd1;
frames[1][6][33] = 8'hd5;
frames[1][6][34] = 8'hd5;
frames[1][6][35] = 8'hd1;
frames[1][6][36] = 8'hd1;
frames[1][6][37] = 8'hd1;
frames[1][6][38] = 8'hd1;
frames[1][6][39] = 8'had;
frames[1][7][0] = 8'hb1;
frames[1][7][1] = 8'hb1;
frames[1][7][2] = 8'hb1;
frames[1][7][3] = 8'hd1;
frames[1][7][4] = 8'hd1;
frames[1][7][5] = 8'hd1;
frames[1][7][6] = 8'hd1;
frames[1][7][7] = 8'hd1;
frames[1][7][8] = 8'hd1;
frames[1][7][9] = 8'hd1;
frames[1][7][10] = 8'hd1;
frames[1][7][11] = 8'hd5;
frames[1][7][12] = 8'hd5;
frames[1][7][13] = 8'hd5;
frames[1][7][14] = 8'hd5;
frames[1][7][15] = 8'hd5;
frames[1][7][16] = 8'hd5;
frames[1][7][17] = 8'hd1;
frames[1][7][18] = 8'h2a;
frames[1][7][19] = 8'h05;
frames[1][7][20] = 8'h05;
frames[1][7][21] = 8'h2a;
frames[1][7][22] = 8'hd1;
frames[1][7][23] = 8'hd5;
frames[1][7][24] = 8'hd5;
frames[1][7][25] = 8'hd5;
frames[1][7][26] = 8'hd5;
frames[1][7][27] = 8'hd5;
frames[1][7][28] = 8'hd1;
frames[1][7][29] = 8'hd1;
frames[1][7][30] = 8'hd1;
frames[1][7][31] = 8'hd1;
frames[1][7][32] = 8'hd1;
frames[1][7][33] = 8'hd5;
frames[1][7][34] = 8'hd5;
frames[1][7][35] = 8'hd5;
frames[1][7][36] = 8'hd1;
frames[1][7][37] = 8'hd1;
frames[1][7][38] = 8'hd1;
frames[1][7][39] = 8'had;
frames[1][8][0] = 8'hb1;
frames[1][8][1] = 8'hb1;
frames[1][8][2] = 8'hd1;
frames[1][8][3] = 8'hd1;
frames[1][8][4] = 8'hd1;
frames[1][8][5] = 8'hd1;
frames[1][8][6] = 8'hd1;
frames[1][8][7] = 8'hd1;
frames[1][8][8] = 8'hd1;
frames[1][8][9] = 8'hd1;
frames[1][8][10] = 8'hd1;
frames[1][8][11] = 8'hd5;
frames[1][8][12] = 8'hd5;
frames[1][8][13] = 8'hd1;
frames[1][8][14] = 8'hd5;
frames[1][8][15] = 8'hf5;
frames[1][8][16] = 8'hd6;
frames[1][8][17] = 8'h8d;
frames[1][8][18] = 8'h05;
frames[1][8][19] = 8'h05;
frames[1][8][20] = 8'h05;
frames[1][8][21] = 8'h06;
frames[1][8][22] = 8'h91;
frames[1][8][23] = 8'hd6;
frames[1][8][24] = 8'hd5;
frames[1][8][25] = 8'hd5;
frames[1][8][26] = 8'hd5;
frames[1][8][27] = 8'hd5;
frames[1][8][28] = 8'hd5;
frames[1][8][29] = 8'hd5;
frames[1][8][30] = 8'hd1;
frames[1][8][31] = 8'hd1;
frames[1][8][32] = 8'hd1;
frames[1][8][33] = 8'hd5;
frames[1][8][34] = 8'hd5;
frames[1][8][35] = 8'hd5;
frames[1][8][36] = 8'hd1;
frames[1][8][37] = 8'hd1;
frames[1][8][38] = 8'hd1;
frames[1][8][39] = 8'had;
frames[1][9][0] = 8'hb1;
frames[1][9][1] = 8'hb1;
frames[1][9][2] = 8'hd1;
frames[1][9][3] = 8'hd1;
frames[1][9][4] = 8'hd1;
frames[1][9][5] = 8'hd1;
frames[1][9][6] = 8'hd1;
frames[1][9][7] = 8'hd1;
frames[1][9][8] = 8'hd1;
frames[1][9][9] = 8'hd1;
frames[1][9][10] = 8'hd1;
frames[1][9][11] = 8'hd5;
frames[1][9][12] = 8'hd5;
frames[1][9][13] = 8'hd1;
frames[1][9][14] = 8'hd5;
frames[1][9][15] = 8'hf5;
frames[1][9][16] = 8'hd6;
frames[1][9][17] = 8'h8d;
frames[1][9][18] = 8'h4e;
frames[1][9][19] = 8'h4e;
frames[1][9][20] = 8'h73;
frames[1][9][21] = 8'h73;
frames[1][9][22] = 8'h91;
frames[1][9][23] = 8'hd6;
frames[1][9][24] = 8'hd5;
frames[1][9][25] = 8'hd5;
frames[1][9][26] = 8'hd5;
frames[1][9][27] = 8'hd5;
frames[1][9][28] = 8'hd5;
frames[1][9][29] = 8'hd5;
frames[1][9][30] = 8'hd1;
frames[1][9][31] = 8'hd1;
frames[1][9][32] = 8'hd1;
frames[1][9][33] = 8'hd5;
frames[1][9][34] = 8'hd5;
frames[1][9][35] = 8'hd5;
frames[1][9][36] = 8'hd1;
frames[1][9][37] = 8'hd1;
frames[1][9][38] = 8'hd1;
frames[1][9][39] = 8'hb1;
frames[1][10][0] = 8'hb1;
frames[1][10][1] = 8'hb1;
frames[1][10][2] = 8'hd1;
frames[1][10][3] = 8'hd1;
frames[1][10][4] = 8'hd1;
frames[1][10][5] = 8'hd1;
frames[1][10][6] = 8'hd1;
frames[1][10][7] = 8'hd1;
frames[1][10][8] = 8'hd1;
frames[1][10][9] = 8'hd1;
frames[1][10][10] = 8'hd1;
frames[1][10][11] = 8'hd5;
frames[1][10][12] = 8'hd1;
frames[1][10][13] = 8'hd1;
frames[1][10][14] = 8'hd5;
frames[1][10][15] = 8'hf5;
frames[1][10][16] = 8'hd6;
frames[1][10][17] = 8'hb1;
frames[1][10][18] = 8'h93;
frames[1][10][19] = 8'h97;
frames[1][10][20] = 8'h73;
frames[1][10][21] = 8'h2a;
frames[1][10][22] = 8'h6d;
frames[1][10][23] = 8'hd6;
frames[1][10][24] = 8'hd5;
frames[1][10][25] = 8'hd5;
frames[1][10][26] = 8'hd5;
frames[1][10][27] = 8'hd5;
frames[1][10][28] = 8'hd5;
frames[1][10][29] = 8'hd5;
frames[1][10][30] = 8'hd1;
frames[1][10][31] = 8'hd1;
frames[1][10][32] = 8'hd1;
frames[1][10][33] = 8'hd1;
frames[1][10][34] = 8'hd5;
frames[1][10][35] = 8'hd5;
frames[1][10][36] = 8'hd1;
frames[1][10][37] = 8'hd1;
frames[1][10][38] = 8'hd1;
frames[1][10][39] = 8'hb1;
frames[1][11][0] = 8'hb1;
frames[1][11][1] = 8'hb1;
frames[1][11][2] = 8'hd1;
frames[1][11][3] = 8'hd1;
frames[1][11][4] = 8'hd1;
frames[1][11][5] = 8'hd1;
frames[1][11][6] = 8'hd1;
frames[1][11][7] = 8'hd1;
frames[1][11][8] = 8'hd1;
frames[1][11][9] = 8'hd1;
frames[1][11][10] = 8'hd1;
frames[1][11][11] = 8'hd5;
frames[1][11][12] = 8'hd1;
frames[1][11][13] = 8'hd1;
frames[1][11][14] = 8'hd5;
frames[1][11][15] = 8'hf5;
frames[1][11][16] = 8'hd6;
frames[1][11][17] = 8'h8d;
frames[1][11][18] = 8'h2a;
frames[1][11][19] = 8'h0a;
frames[1][11][20] = 8'h05;
frames[1][11][21] = 8'h05;
frames[1][11][22] = 8'h8d;
frames[1][11][23] = 8'hd6;
frames[1][11][24] = 8'hd5;
frames[1][11][25] = 8'hd5;
frames[1][11][26] = 8'hd5;
frames[1][11][27] = 8'hd5;
frames[1][11][28] = 8'hd5;
frames[1][11][29] = 8'hd5;
frames[1][11][30] = 8'hd1;
frames[1][11][31] = 8'hd1;
frames[1][11][32] = 8'hd1;
frames[1][11][33] = 8'hd1;
frames[1][11][34] = 8'hd5;
frames[1][11][35] = 8'hd5;
frames[1][11][36] = 8'hd1;
frames[1][11][37] = 8'hd1;
frames[1][11][38] = 8'hd1;
frames[1][11][39] = 8'hb1;
frames[1][12][0] = 8'had;
frames[1][12][1] = 8'hb1;
frames[1][12][2] = 8'hd1;
frames[1][12][3] = 8'hd1;
frames[1][12][4] = 8'hd1;
frames[1][12][5] = 8'hd1;
frames[1][12][6] = 8'hd1;
frames[1][12][7] = 8'hd1;
frames[1][12][8] = 8'hd1;
frames[1][12][9] = 8'hd1;
frames[1][12][10] = 8'hd1;
frames[1][12][11] = 8'hd5;
frames[1][12][12] = 8'hd1;
frames[1][12][13] = 8'hd1;
frames[1][12][14] = 8'hd5;
frames[1][12][15] = 8'hd5;
frames[1][12][16] = 8'hd5;
frames[1][12][17] = 8'hd1;
frames[1][12][18] = 8'h2a;
frames[1][12][19] = 8'h05;
frames[1][12][20] = 8'h05;
frames[1][12][21] = 8'h2a;
frames[1][12][22] = 8'hd5;
frames[1][12][23] = 8'hd5;
frames[1][12][24] = 8'hd5;
frames[1][12][25] = 8'hd5;
frames[1][12][26] = 8'hf5;
frames[1][12][27] = 8'hd5;
frames[1][12][28] = 8'hd5;
frames[1][12][29] = 8'hd1;
frames[1][12][30] = 8'hd1;
frames[1][12][31] = 8'hd1;
frames[1][12][32] = 8'hd1;
frames[1][12][33] = 8'hd1;
frames[1][12][34] = 8'hd5;
frames[1][12][35] = 8'hd5;
frames[1][12][36] = 8'hd1;
frames[1][12][37] = 8'hd1;
frames[1][12][38] = 8'hd1;
frames[1][12][39] = 8'hb1;
frames[1][13][0] = 8'had;
frames[1][13][1] = 8'hb1;
frames[1][13][2] = 8'hd1;
frames[1][13][3] = 8'hd1;
frames[1][13][4] = 8'hd1;
frames[1][13][5] = 8'hd1;
frames[1][13][6] = 8'hd1;
frames[1][13][7] = 8'hd1;
frames[1][13][8] = 8'hd1;
frames[1][13][9] = 8'hd1;
frames[1][13][10] = 8'hd1;
frames[1][13][11] = 8'hd5;
frames[1][13][12] = 8'hd1;
frames[1][13][13] = 8'hd1;
frames[1][13][14] = 8'hd5;
frames[1][13][15] = 8'hd5;
frames[1][13][16] = 8'hd5;
frames[1][13][17] = 8'hd5;
frames[1][13][18] = 8'hb2;
frames[1][13][19] = 8'h6d;
frames[1][13][20] = 8'h6d;
frames[1][13][21] = 8'h91;
frames[1][13][22] = 8'hd5;
frames[1][13][23] = 8'hd5;
frames[1][13][24] = 8'hd5;
frames[1][13][25] = 8'hd5;
frames[1][13][26] = 8'hd5;
frames[1][13][27] = 8'hd5;
frames[1][13][28] = 8'hd5;
frames[1][13][29] = 8'hd5;
frames[1][13][30] = 8'hd1;
frames[1][13][31] = 8'hd1;
frames[1][13][32] = 8'hd1;
frames[1][13][33] = 8'hd1;
frames[1][13][34] = 8'hd5;
frames[1][13][35] = 8'hd5;
frames[1][13][36] = 8'hd1;
frames[1][13][37] = 8'hd1;
frames[1][13][38] = 8'hb1;
frames[1][13][39] = 8'hb1;
frames[1][14][0] = 8'had;
frames[1][14][1] = 8'hb1;
frames[1][14][2] = 8'hd1;
frames[1][14][3] = 8'hd1;
frames[1][14][4] = 8'hd1;
frames[1][14][5] = 8'hd1;
frames[1][14][6] = 8'hd1;
frames[1][14][7] = 8'hd1;
frames[1][14][8] = 8'hd1;
frames[1][14][9] = 8'hd1;
frames[1][14][10] = 8'hd1;
frames[1][14][11] = 8'hd1;
frames[1][14][12] = 8'hd5;
frames[1][14][13] = 8'hd5;
frames[1][14][14] = 8'hd5;
frames[1][14][15] = 8'hd5;
frames[1][14][16] = 8'hf5;
frames[1][14][17] = 8'hd5;
frames[1][14][18] = 8'hfa;
frames[1][14][19] = 8'hfa;
frames[1][14][20] = 8'hf5;
frames[1][14][21] = 8'hf5;
frames[1][14][22] = 8'hfa;
frames[1][14][23] = 8'hfa;
frames[1][14][24] = 8'hf5;
frames[1][14][25] = 8'hd5;
frames[1][14][26] = 8'hd5;
frames[1][14][27] = 8'hd5;
frames[1][14][28] = 8'hd5;
frames[1][14][29] = 8'hd5;
frames[1][14][30] = 8'hd1;
frames[1][14][31] = 8'hd1;
frames[1][14][32] = 8'hd1;
frames[1][14][33] = 8'hd1;
frames[1][14][34] = 8'hd1;
frames[1][14][35] = 8'hd5;
frames[1][14][36] = 8'hd1;
frames[1][14][37] = 8'hd1;
frames[1][14][38] = 8'hb1;
frames[1][14][39] = 8'hb1;
frames[1][15][0] = 8'had;
frames[1][15][1] = 8'hb1;
frames[1][15][2] = 8'hd1;
frames[1][15][3] = 8'hd1;
frames[1][15][4] = 8'hd1;
frames[1][15][5] = 8'hd1;
frames[1][15][6] = 8'hd1;
frames[1][15][7] = 8'hd1;
frames[1][15][8] = 8'hd1;
frames[1][15][9] = 8'hd1;
frames[1][15][10] = 8'hd1;
frames[1][15][11] = 8'hd1;
frames[1][15][12] = 8'hd5;
frames[1][15][13] = 8'hd5;
frames[1][15][14] = 8'hd5;
frames[1][15][15] = 8'hd5;
frames[1][15][16] = 8'hf6;
frames[1][15][17] = 8'hf6;
frames[1][15][18] = 8'hfa;
frames[1][15][19] = 8'hfa;
frames[1][15][20] = 8'hf6;
frames[1][15][21] = 8'hfa;
frames[1][15][22] = 8'hfa;
frames[1][15][23] = 8'hfa;
frames[1][15][24] = 8'hd5;
frames[1][15][25] = 8'hd5;
frames[1][15][26] = 8'hd5;
frames[1][15][27] = 8'hd5;
frames[1][15][28] = 8'hd5;
frames[1][15][29] = 8'hd5;
frames[1][15][30] = 8'hd1;
frames[1][15][31] = 8'hd1;
frames[1][15][32] = 8'hd1;
frames[1][15][33] = 8'hd1;
frames[1][15][34] = 8'hd1;
frames[1][15][35] = 8'hd1;
frames[1][15][36] = 8'hd1;
frames[1][15][37] = 8'hd1;
frames[1][15][38] = 8'hb1;
frames[1][15][39] = 8'hb1;
frames[1][16][0] = 8'had;
frames[1][16][1] = 8'hb1;
frames[1][16][2] = 8'hb1;
frames[1][16][3] = 8'hb1;
frames[1][16][4] = 8'hd1;
frames[1][16][5] = 8'hd1;
frames[1][16][6] = 8'hd1;
frames[1][16][7] = 8'hd1;
frames[1][16][8] = 8'hd1;
frames[1][16][9] = 8'hd1;
frames[1][16][10] = 8'hd5;
frames[1][16][11] = 8'hd5;
frames[1][16][12] = 8'hd1;
frames[1][16][13] = 8'hd1;
frames[1][16][14] = 8'hd5;
frames[1][16][15] = 8'hf5;
frames[1][16][16] = 8'hd5;
frames[1][16][17] = 8'hd5;
frames[1][16][18] = 8'hd5;
frames[1][16][19] = 8'hf6;
frames[1][16][20] = 8'hd5;
frames[1][16][21] = 8'hd5;
frames[1][16][22] = 8'hf6;
frames[1][16][23] = 8'hf6;
frames[1][16][24] = 8'hf5;
frames[1][16][25] = 8'hd5;
frames[1][16][26] = 8'hd5;
frames[1][16][27] = 8'hd5;
frames[1][16][28] = 8'hd5;
frames[1][16][29] = 8'hd5;
frames[1][16][30] = 8'hd1;
frames[1][16][31] = 8'hd1;
frames[1][16][32] = 8'hd1;
frames[1][16][33] = 8'hd1;
frames[1][16][34] = 8'hd1;
frames[1][16][35] = 8'hd1;
frames[1][16][36] = 8'hd1;
frames[1][16][37] = 8'hb1;
frames[1][16][38] = 8'hb1;
frames[1][16][39] = 8'hb1;
frames[1][17][0] = 8'had;
frames[1][17][1] = 8'hb1;
frames[1][17][2] = 8'hb1;
frames[1][17][3] = 8'hb1;
frames[1][17][4] = 8'hd1;
frames[1][17][5] = 8'hd1;
frames[1][17][6] = 8'hd1;
frames[1][17][7] = 8'hd1;
frames[1][17][8] = 8'hd1;
frames[1][17][9] = 8'hd1;
frames[1][17][10] = 8'hd5;
frames[1][17][11] = 8'hd5;
frames[1][17][12] = 8'hd1;
frames[1][17][13] = 8'hd1;
frames[1][17][14] = 8'hd6;
frames[1][17][15] = 8'hfa;
frames[1][17][16] = 8'hfa;
frames[1][17][17] = 8'hd6;
frames[1][17][18] = 8'hf6;
frames[1][17][19] = 8'hfa;
frames[1][17][20] = 8'hd6;
frames[1][17][21] = 8'hf6;
frames[1][17][22] = 8'hfa;
frames[1][17][23] = 8'hfa;
frames[1][17][24] = 8'hfa;
frames[1][17][25] = 8'hd6;
frames[1][17][26] = 8'hd5;
frames[1][17][27] = 8'hd5;
frames[1][17][28] = 8'hd5;
frames[1][17][29] = 8'hd5;
frames[1][17][30] = 8'hd1;
frames[1][17][31] = 8'hd1;
frames[1][17][32] = 8'hd1;
frames[1][17][33] = 8'hd1;
frames[1][17][34] = 8'hd1;
frames[1][17][35] = 8'hd1;
frames[1][17][36] = 8'hd1;
frames[1][17][37] = 8'hb1;
frames[1][17][38] = 8'hb1;
frames[1][17][39] = 8'hb1;
frames[1][18][0] = 8'had;
frames[1][18][1] = 8'hb1;
frames[1][18][2] = 8'hb1;
frames[1][18][3] = 8'hb1;
frames[1][18][4] = 8'hd1;
frames[1][18][5] = 8'hd1;
frames[1][18][6] = 8'hd1;
frames[1][18][7] = 8'hd1;
frames[1][18][8] = 8'hd1;
frames[1][18][9] = 8'hd1;
frames[1][18][10] = 8'hd5;
frames[1][18][11] = 8'hd5;
frames[1][18][12] = 8'hd5;
frames[1][18][13] = 8'hd1;
frames[1][18][14] = 8'hd6;
frames[1][18][15] = 8'hfa;
frames[1][18][16] = 8'hfa;
frames[1][18][17] = 8'hd6;
frames[1][18][18] = 8'hf6;
frames[1][18][19] = 8'hfa;
frames[1][18][20] = 8'hd6;
frames[1][18][21] = 8'hfa;
frames[1][18][22] = 8'hfa;
frames[1][18][23] = 8'hda;
frames[1][18][24] = 8'hfa;
frames[1][18][25] = 8'hf6;
frames[1][18][26] = 8'hd5;
frames[1][18][27] = 8'hd5;
frames[1][18][28] = 8'hd5;
frames[1][18][29] = 8'hd1;
frames[1][18][30] = 8'hd1;
frames[1][18][31] = 8'hd1;
frames[1][18][32] = 8'hd1;
frames[1][18][33] = 8'hd1;
frames[1][18][34] = 8'hd1;
frames[1][18][35] = 8'hd1;
frames[1][18][36] = 8'hd1;
frames[1][18][37] = 8'hb1;
frames[1][18][38] = 8'hb1;
frames[1][18][39] = 8'hb1;
frames[1][19][0] = 8'hac;
frames[1][19][1] = 8'hb1;
frames[1][19][2] = 8'hb1;
frames[1][19][3] = 8'hb1;
frames[1][19][4] = 8'hd1;
frames[1][19][5] = 8'hd1;
frames[1][19][6] = 8'hd1;
frames[1][19][7] = 8'hd1;
frames[1][19][8] = 8'hd1;
frames[1][19][9] = 8'hd1;
frames[1][19][10] = 8'hd5;
frames[1][19][11] = 8'hd5;
frames[1][19][12] = 8'hd5;
frames[1][19][13] = 8'hd1;
frames[1][19][14] = 8'hd6;
frames[1][19][15] = 8'hfa;
frames[1][19][16] = 8'hfa;
frames[1][19][17] = 8'hda;
frames[1][19][18] = 8'hfa;
frames[1][19][19] = 8'hfa;
frames[1][19][20] = 8'hd5;
frames[1][19][21] = 8'hd5;
frames[1][19][22] = 8'hfa;
frames[1][19][23] = 8'hfa;
frames[1][19][24] = 8'hfa;
frames[1][19][25] = 8'hd6;
frames[1][19][26] = 8'hd5;
frames[1][19][27] = 8'hd5;
frames[1][19][28] = 8'hd1;
frames[1][19][29] = 8'hd1;
frames[1][19][30] = 8'hd1;
frames[1][19][31] = 8'hd1;
frames[1][19][32] = 8'hd1;
frames[1][19][33] = 8'hd1;
frames[1][19][34] = 8'hd1;
frames[1][19][35] = 8'hd1;
frames[1][19][36] = 8'hd1;
frames[1][19][37] = 8'hb1;
frames[1][19][38] = 8'hb1;
frames[1][19][39] = 8'hb1;
frames[1][20][0] = 8'hac;
frames[1][20][1] = 8'hb1;
frames[1][20][2] = 8'hb1;
frames[1][20][3] = 8'hb1;
frames[1][20][4] = 8'hd1;
frames[1][20][5] = 8'hd1;
frames[1][20][6] = 8'hd1;
frames[1][20][7] = 8'hd1;
frames[1][20][8] = 8'hd1;
frames[1][20][9] = 8'hd1;
frames[1][20][10] = 8'hd5;
frames[1][20][11] = 8'hd5;
frames[1][20][12] = 8'hd5;
frames[1][20][13] = 8'hd5;
frames[1][20][14] = 8'hd5;
frames[1][20][15] = 8'hf5;
frames[1][20][16] = 8'hd6;
frames[1][20][17] = 8'hf6;
frames[1][20][18] = 8'hf6;
frames[1][20][19] = 8'hf6;
frames[1][20][20] = 8'hd5;
frames[1][20][21] = 8'hd5;
frames[1][20][22] = 8'hd6;
frames[1][20][23] = 8'hf6;
frames[1][20][24] = 8'hf6;
frames[1][20][25] = 8'hd5;
frames[1][20][26] = 8'hd5;
frames[1][20][27] = 8'hd5;
frames[1][20][28] = 8'hd5;
frames[1][20][29] = 8'hd1;
frames[1][20][30] = 8'hd1;
frames[1][20][31] = 8'hd1;
frames[1][20][32] = 8'hd1;
frames[1][20][33] = 8'hd1;
frames[1][20][34] = 8'hd1;
frames[1][20][35] = 8'hd1;
frames[1][20][36] = 8'hb1;
frames[1][20][37] = 8'hb1;
frames[1][20][38] = 8'hb1;
frames[1][20][39] = 8'hb1;
frames[1][21][0] = 8'hac;
frames[1][21][1] = 8'hb1;
frames[1][21][2] = 8'hb1;
frames[1][21][3] = 8'hb1;
frames[1][21][4] = 8'hd1;
frames[1][21][5] = 8'hd1;
frames[1][21][6] = 8'hd1;
frames[1][21][7] = 8'hd1;
frames[1][21][8] = 8'hd1;
frames[1][21][9] = 8'hd1;
frames[1][21][10] = 8'hd1;
frames[1][21][11] = 8'hd1;
frames[1][21][12] = 8'hd5;
frames[1][21][13] = 8'hd5;
frames[1][21][14] = 8'hd5;
frames[1][21][15] = 8'hfa;
frames[1][21][16] = 8'hfa;
frames[1][21][17] = 8'hfa;
frames[1][21][18] = 8'hfa;
frames[1][21][19] = 8'hfa;
frames[1][21][20] = 8'hfa;
frames[1][21][21] = 8'hf6;
frames[1][21][22] = 8'hd6;
frames[1][21][23] = 8'hfa;
frames[1][21][24] = 8'hf6;
frames[1][21][25] = 8'hd5;
frames[1][21][26] = 8'hd5;
frames[1][21][27] = 8'hd5;
frames[1][21][28] = 8'hd5;
frames[1][21][29] = 8'hd1;
frames[1][21][30] = 8'hd1;
frames[1][21][31] = 8'hd1;
frames[1][21][32] = 8'hd1;
frames[1][21][33] = 8'hd1;
frames[1][21][34] = 8'hb1;
frames[1][21][35] = 8'hd1;
frames[1][21][36] = 8'hb1;
frames[1][21][37] = 8'hb1;
frames[1][21][38] = 8'hb1;
frames[1][21][39] = 8'hb1;
frames[1][22][0] = 8'hac;
frames[1][22][1] = 8'hb1;
frames[1][22][2] = 8'hb1;
frames[1][22][3] = 8'hb1;
frames[1][22][4] = 8'hb1;
frames[1][22][5] = 8'hd1;
frames[1][22][6] = 8'hd1;
frames[1][22][7] = 8'hd1;
frames[1][22][8] = 8'hd1;
frames[1][22][9] = 8'hd1;
frames[1][22][10] = 8'hd1;
frames[1][22][11] = 8'hd1;
frames[1][22][12] = 8'hd1;
frames[1][22][13] = 8'hd5;
frames[1][22][14] = 8'hd5;
frames[1][22][15] = 8'hfa;
frames[1][22][16] = 8'hfa;
frames[1][22][17] = 8'hda;
frames[1][22][18] = 8'hd6;
frames[1][22][19] = 8'hfa;
frames[1][22][20] = 8'hfa;
frames[1][22][21] = 8'hfa;
frames[1][22][22] = 8'hd6;
frames[1][22][23] = 8'hfa;
frames[1][22][24] = 8'hf6;
frames[1][22][25] = 8'hd5;
frames[1][22][26] = 8'hd5;
frames[1][22][27] = 8'hd1;
frames[1][22][28] = 8'hd1;
frames[1][22][29] = 8'hd1;
frames[1][22][30] = 8'hd1;
frames[1][22][31] = 8'hd1;
frames[1][22][32] = 8'hd1;
frames[1][22][33] = 8'hd1;
frames[1][22][34] = 8'hb1;
frames[1][22][35] = 8'hd1;
frames[1][22][36] = 8'hb1;
frames[1][22][37] = 8'hb1;
frames[1][22][38] = 8'hb1;
frames[1][22][39] = 8'hb1;
frames[1][23][0] = 8'hac;
frames[1][23][1] = 8'hb1;
frames[1][23][2] = 8'hb1;
frames[1][23][3] = 8'hb1;
frames[1][23][4] = 8'hb1;
frames[1][23][5] = 8'hd1;
frames[1][23][6] = 8'hd1;
frames[1][23][7] = 8'hd1;
frames[1][23][8] = 8'hd1;
frames[1][23][9] = 8'hd1;
frames[1][23][10] = 8'hd1;
frames[1][23][11] = 8'hd1;
frames[1][23][12] = 8'hd1;
frames[1][23][13] = 8'hd5;
frames[1][23][14] = 8'hd5;
frames[1][23][15] = 8'hfa;
frames[1][23][16] = 8'hfa;
frames[1][23][17] = 8'hfa;
frames[1][23][18] = 8'hfa;
frames[1][23][19] = 8'hfa;
frames[1][23][20] = 8'hfa;
frames[1][23][21] = 8'hfa;
frames[1][23][22] = 8'hfa;
frames[1][23][23] = 8'hfa;
frames[1][23][24] = 8'hfa;
frames[1][23][25] = 8'hd5;
frames[1][23][26] = 8'hd1;
frames[1][23][27] = 8'hd1;
frames[1][23][28] = 8'hd1;
frames[1][23][29] = 8'hd1;
frames[1][23][30] = 8'hd1;
frames[1][23][31] = 8'hd1;
frames[1][23][32] = 8'hd1;
frames[1][23][33] = 8'hb1;
frames[1][23][34] = 8'hb1;
frames[1][23][35] = 8'hd1;
frames[1][23][36] = 8'hb1;
frames[1][23][37] = 8'hb1;
frames[1][23][38] = 8'hb1;
frames[1][23][39] = 8'hb1;
frames[1][24][0] = 8'hac;
frames[1][24][1] = 8'hb1;
frames[1][24][2] = 8'hb1;
frames[1][24][3] = 8'hb1;
frames[1][24][4] = 8'hb1;
frames[1][24][5] = 8'hd1;
frames[1][24][6] = 8'hd1;
frames[1][24][7] = 8'hd1;
frames[1][24][8] = 8'hd1;
frames[1][24][9] = 8'hd1;
frames[1][24][10] = 8'hd1;
frames[1][24][11] = 8'hd1;
frames[1][24][12] = 8'hd1;
frames[1][24][13] = 8'hd1;
frames[1][24][14] = 8'hd5;
frames[1][24][15] = 8'hd5;
frames[1][24][16] = 8'hd5;
frames[1][24][17] = 8'hd5;
frames[1][24][18] = 8'hd5;
frames[1][24][19] = 8'hd5;
frames[1][24][20] = 8'hd5;
frames[1][24][21] = 8'hd5;
frames[1][24][22] = 8'hd5;
frames[1][24][23] = 8'hd5;
frames[1][24][24] = 8'hd5;
frames[1][24][25] = 8'hd5;
frames[1][24][26] = 8'hd1;
frames[1][24][27] = 8'hd1;
frames[1][24][28] = 8'hd1;
frames[1][24][29] = 8'hd1;
frames[1][24][30] = 8'hd1;
frames[1][24][31] = 8'hd1;
frames[1][24][32] = 8'hb1;
frames[1][24][33] = 8'hb1;
frames[1][24][34] = 8'hb1;
frames[1][24][35] = 8'hd1;
frames[1][24][36] = 8'hb1;
frames[1][24][37] = 8'hb1;
frames[1][24][38] = 8'hb1;
frames[1][24][39] = 8'hb1;
frames[1][25][0] = 8'hac;
frames[1][25][1] = 8'hac;
frames[1][25][2] = 8'hac;
frames[1][25][3] = 8'hac;
frames[1][25][4] = 8'hb1;
frames[1][25][5] = 8'hd1;
frames[1][25][6] = 8'hd1;
frames[1][25][7] = 8'hd1;
frames[1][25][8] = 8'hd1;
frames[1][25][9] = 8'hd1;
frames[1][25][10] = 8'hd1;
frames[1][25][11] = 8'hd1;
frames[1][25][12] = 8'hd1;
frames[1][25][13] = 8'hd1;
frames[1][25][14] = 8'hd1;
frames[1][25][15] = 8'hd1;
frames[1][25][16] = 8'hd1;
frames[1][25][17] = 8'hd1;
frames[1][25][18] = 8'hd1;
frames[1][25][19] = 8'hd5;
frames[1][25][20] = 8'hd5;
frames[1][25][21] = 8'hd5;
frames[1][25][22] = 8'hd5;
frames[1][25][23] = 8'hd5;
frames[1][25][24] = 8'hd5;
frames[1][25][25] = 8'hd5;
frames[1][25][26] = 8'hd1;
frames[1][25][27] = 8'hd1;
frames[1][25][28] = 8'hd1;
frames[1][25][29] = 8'hd1;
frames[1][25][30] = 8'hd1;
frames[1][25][31] = 8'hd1;
frames[1][25][32] = 8'hb1;
frames[1][25][33] = 8'hb1;
frames[1][25][34] = 8'hb1;
frames[1][25][35] = 8'hb1;
frames[1][25][36] = 8'hb1;
frames[1][25][37] = 8'hb1;
frames[1][25][38] = 8'hb1;
frames[1][25][39] = 8'hb1;
frames[1][26][0] = 8'h8c;
frames[1][26][1] = 8'hac;
frames[1][26][2] = 8'hac;
frames[1][26][3] = 8'hac;
frames[1][26][4] = 8'hb0;
frames[1][26][5] = 8'hb1;
frames[1][26][6] = 8'hd1;
frames[1][26][7] = 8'hd1;
frames[1][26][8] = 8'hd1;
frames[1][26][9] = 8'hd1;
frames[1][26][10] = 8'hd1;
frames[1][26][11] = 8'hd1;
frames[1][26][12] = 8'hd1;
frames[1][26][13] = 8'hd1;
frames[1][26][14] = 8'hd1;
frames[1][26][15] = 8'hd1;
frames[1][26][16] = 8'hd1;
frames[1][26][17] = 8'hd1;
frames[1][26][18] = 8'hd1;
frames[1][26][19] = 8'hd1;
frames[1][26][20] = 8'hd1;
frames[1][26][21] = 8'hd1;
frames[1][26][22] = 8'hd5;
frames[1][26][23] = 8'hd5;
frames[1][26][24] = 8'hd5;
frames[1][26][25] = 8'hd1;
frames[1][26][26] = 8'hd1;
frames[1][26][27] = 8'hd1;
frames[1][26][28] = 8'hd1;
frames[1][26][29] = 8'hd1;
frames[1][26][30] = 8'hd1;
frames[1][26][31] = 8'hb1;
frames[1][26][32] = 8'hb1;
frames[1][26][33] = 8'hb1;
frames[1][26][34] = 8'hb1;
frames[1][26][35] = 8'hb1;
frames[1][26][36] = 8'hb1;
frames[1][26][37] = 8'hb1;
frames[1][26][38] = 8'hb1;
frames[1][26][39] = 8'hb1;
frames[1][27][0] = 8'h8c;
frames[1][27][1] = 8'hac;
frames[1][27][2] = 8'hac;
frames[1][27][3] = 8'hac;
frames[1][27][4] = 8'hac;
frames[1][27][5] = 8'hb1;
frames[1][27][6] = 8'hd1;
frames[1][27][7] = 8'hd1;
frames[1][27][8] = 8'hd1;
frames[1][27][9] = 8'hd1;
frames[1][27][10] = 8'hd1;
frames[1][27][11] = 8'hd1;
frames[1][27][12] = 8'hd1;
frames[1][27][13] = 8'hd1;
frames[1][27][14] = 8'hd1;
frames[1][27][15] = 8'hd1;
frames[1][27][16] = 8'hb1;
frames[1][27][17] = 8'hb1;
frames[1][27][18] = 8'hb1;
frames[1][27][19] = 8'hd1;
frames[1][27][20] = 8'hd1;
frames[1][27][21] = 8'hd1;
frames[1][27][22] = 8'hd1;
frames[1][27][23] = 8'hd1;
frames[1][27][24] = 8'hd1;
frames[1][27][25] = 8'hd1;
frames[1][27][26] = 8'hd1;
frames[1][27][27] = 8'hd1;
frames[1][27][28] = 8'hd1;
frames[1][27][29] = 8'hd1;
frames[1][27][30] = 8'hd1;
frames[1][27][31] = 8'hb1;
frames[1][27][32] = 8'hb1;
frames[1][27][33] = 8'hb1;
frames[1][27][34] = 8'hb1;
frames[1][27][35] = 8'hb1;
frames[1][27][36] = 8'hb1;
frames[1][27][37] = 8'hb1;
frames[1][27][38] = 8'hb1;
frames[1][27][39] = 8'hb1;
frames[1][28][0] = 8'h8c;
frames[1][28][1] = 8'h8c;
frames[1][28][2] = 8'h8c;
frames[1][28][3] = 8'hac;
frames[1][28][4] = 8'hac;
frames[1][28][5] = 8'had;
frames[1][28][6] = 8'hb1;
frames[1][28][7] = 8'hb1;
frames[1][28][8] = 8'hd1;
frames[1][28][9] = 8'hd1;
frames[1][28][10] = 8'hd1;
frames[1][28][11] = 8'hd1;
frames[1][28][12] = 8'hd1;
frames[1][28][13] = 8'hd1;
frames[1][28][14] = 8'hd1;
frames[1][28][15] = 8'hd1;
frames[1][28][16] = 8'had;
frames[1][28][17] = 8'hac;
frames[1][28][18] = 8'had;
frames[1][28][19] = 8'had;
frames[1][28][20] = 8'hb1;
frames[1][28][21] = 8'hb1;
frames[1][28][22] = 8'hd1;
frames[1][28][23] = 8'hd1;
frames[1][28][24] = 8'hd1;
frames[1][28][25] = 8'hd1;
frames[1][28][26] = 8'hd1;
frames[1][28][27] = 8'hb1;
frames[1][28][28] = 8'hb1;
frames[1][28][29] = 8'hb1;
frames[1][28][30] = 8'hb1;
frames[1][28][31] = 8'hb1;
frames[1][28][32] = 8'hb1;
frames[1][28][33] = 8'hb1;
frames[1][28][34] = 8'hb1;
frames[1][28][35] = 8'hb1;
frames[1][28][36] = 8'hb1;
frames[1][28][37] = 8'hb1;
frames[1][28][38] = 8'hb1;
frames[1][28][39] = 8'had;
frames[1][29][0] = 8'h8c;
frames[1][29][1] = 8'h8c;
frames[1][29][2] = 8'h8c;
frames[1][29][3] = 8'h8c;
frames[1][29][4] = 8'hac;
frames[1][29][5] = 8'hac;
frames[1][29][6] = 8'hac;
frames[1][29][7] = 8'hb1;
frames[1][29][8] = 8'hd1;
frames[1][29][9] = 8'hd1;
frames[1][29][10] = 8'hd1;
frames[1][29][11] = 8'hd1;
frames[1][29][12] = 8'hd1;
frames[1][29][13] = 8'hd1;
frames[1][29][14] = 8'hd1;
frames[1][29][15] = 8'hd1;
frames[1][29][16] = 8'had;
frames[1][29][17] = 8'hac;
frames[1][29][18] = 8'hac;
frames[1][29][19] = 8'hac;
frames[1][29][20] = 8'hac;
frames[1][29][21] = 8'hac;
frames[1][29][22] = 8'hb1;
frames[1][29][23] = 8'hd1;
frames[1][29][24] = 8'hd1;
frames[1][29][25] = 8'hd1;
frames[1][29][26] = 8'hb1;
frames[1][29][27] = 8'hb1;
frames[1][29][28] = 8'hb1;
frames[1][29][29] = 8'hb1;
frames[1][29][30] = 8'hb1;
frames[1][29][31] = 8'hb1;
frames[1][29][32] = 8'hb1;
frames[1][29][33] = 8'hb1;
frames[1][29][34] = 8'hb1;
frames[1][29][35] = 8'hb1;
frames[1][29][36] = 8'hb1;
frames[1][29][37] = 8'hb1;
frames[1][29][38] = 8'hb1;
frames[1][29][39] = 8'hb1;
frames[2][0][0] = 8'hd1;
frames[2][0][1] = 8'hb1;
frames[2][0][2] = 8'hb1;
frames[2][0][3] = 8'hd1;
frames[2][0][4] = 8'hd1;
frames[2][0][5] = 8'hd1;
frames[2][0][6] = 8'hd5;
frames[2][0][7] = 8'hd5;
frames[2][0][8] = 8'hd5;
frames[2][0][9] = 8'hd1;
frames[2][0][10] = 8'hd1;
frames[2][0][11] = 8'hd5;
frames[2][0][12] = 8'hd5;
frames[2][0][13] = 8'hd5;
frames[2][0][14] = 8'hd5;
frames[2][0][15] = 8'hd5;
frames[2][0][16] = 8'hd5;
frames[2][0][17] = 8'hd1;
frames[2][0][18] = 8'hd5;
frames[2][0][19] = 8'hd1;
frames[2][0][20] = 8'hd1;
frames[2][0][21] = 8'hd1;
frames[2][0][22] = 8'hd5;
frames[2][0][23] = 8'hd5;
frames[2][0][24] = 8'hd5;
frames[2][0][25] = 8'hd5;
frames[2][0][26] = 8'hd1;
frames[2][0][27] = 8'hd1;
frames[2][0][28] = 8'hd1;
frames[2][0][29] = 8'hd1;
frames[2][0][30] = 8'hd1;
frames[2][0][31] = 8'hd1;
frames[2][0][32] = 8'hd1;
frames[2][0][33] = 8'hd5;
frames[2][0][34] = 8'hd5;
frames[2][0][35] = 8'hd1;
frames[2][0][36] = 8'hd1;
frames[2][0][37] = 8'hd1;
frames[2][0][38] = 8'hb1;
frames[2][0][39] = 8'had;
frames[2][1][0] = 8'had;
frames[2][1][1] = 8'hd1;
frames[2][1][2] = 8'hd1;
frames[2][1][3] = 8'hb1;
frames[2][1][4] = 8'hb1;
frames[2][1][5] = 8'hd1;
frames[2][1][6] = 8'hd1;
frames[2][1][7] = 8'hd5;
frames[2][1][8] = 8'hd1;
frames[2][1][9] = 8'hd1;
frames[2][1][10] = 8'hd1;
frames[2][1][11] = 8'hd5;
frames[2][1][12] = 8'hd5;
frames[2][1][13] = 8'hd5;
frames[2][1][14] = 8'hd5;
frames[2][1][15] = 8'hd5;
frames[2][1][16] = 8'hd5;
frames[2][1][17] = 8'hd1;
frames[2][1][18] = 8'hd1;
frames[2][1][19] = 8'hd1;
frames[2][1][20] = 8'hd1;
frames[2][1][21] = 8'hd1;
frames[2][1][22] = 8'hd5;
frames[2][1][23] = 8'hd5;
frames[2][1][24] = 8'hd5;
frames[2][1][25] = 8'hd5;
frames[2][1][26] = 8'hd1;
frames[2][1][27] = 8'hd1;
frames[2][1][28] = 8'hd1;
frames[2][1][29] = 8'hd1;
frames[2][1][30] = 8'hd1;
frames[2][1][31] = 8'hd1;
frames[2][1][32] = 8'hd1;
frames[2][1][33] = 8'hd5;
frames[2][1][34] = 8'hd5;
frames[2][1][35] = 8'hd1;
frames[2][1][36] = 8'hd1;
frames[2][1][37] = 8'hd1;
frames[2][1][38] = 8'hb1;
frames[2][1][39] = 8'had;
frames[2][2][0] = 8'h8d;
frames[2][2][1] = 8'had;
frames[2][2][2] = 8'hd1;
frames[2][2][3] = 8'hd1;
frames[2][2][4] = 8'hd1;
frames[2][2][5] = 8'hd5;
frames[2][2][6] = 8'hf6;
frames[2][2][7] = 8'hd6;
frames[2][2][8] = 8'hd1;
frames[2][2][9] = 8'hd1;
frames[2][2][10] = 8'hd1;
frames[2][2][11] = 8'hd5;
frames[2][2][12] = 8'hd5;
frames[2][2][13] = 8'hd5;
frames[2][2][14] = 8'hd5;
frames[2][2][15] = 8'hd5;
frames[2][2][16] = 8'hd1;
frames[2][2][17] = 8'hd1;
frames[2][2][18] = 8'hd1;
frames[2][2][19] = 8'hd1;
frames[2][2][20] = 8'hd1;
frames[2][2][21] = 8'hd1;
frames[2][2][22] = 8'hd5;
frames[2][2][23] = 8'hd5;
frames[2][2][24] = 8'hd5;
frames[2][2][25] = 8'hd5;
frames[2][2][26] = 8'hd5;
frames[2][2][27] = 8'hd1;
frames[2][2][28] = 8'hd1;
frames[2][2][29] = 8'hd1;
frames[2][2][30] = 8'hd1;
frames[2][2][31] = 8'hd1;
frames[2][2][32] = 8'hd1;
frames[2][2][33] = 8'hd5;
frames[2][2][34] = 8'hd1;
frames[2][2][35] = 8'hd1;
frames[2][2][36] = 8'hd1;
frames[2][2][37] = 8'hd1;
frames[2][2][38] = 8'hb1;
frames[2][2][39] = 8'had;
frames[2][3][0] = 8'h8d;
frames[2][3][1] = 8'h89;
frames[2][3][2] = 8'h8d;
frames[2][3][3] = 8'had;
frames[2][3][4] = 8'hb1;
frames[2][3][5] = 8'hb1;
frames[2][3][6] = 8'had;
frames[2][3][7] = 8'had;
frames[2][3][8] = 8'hd1;
frames[2][3][9] = 8'hd1;
frames[2][3][10] = 8'hd1;
frames[2][3][11] = 8'hd5;
frames[2][3][12] = 8'hd5;
frames[2][3][13] = 8'hd5;
frames[2][3][14] = 8'hd5;
frames[2][3][15] = 8'hd5;
frames[2][3][16] = 8'hd1;
frames[2][3][17] = 8'hd1;
frames[2][3][18] = 8'hd1;
frames[2][3][19] = 8'hd1;
frames[2][3][20] = 8'hd1;
frames[2][3][21] = 8'hd1;
frames[2][3][22] = 8'hd5;
frames[2][3][23] = 8'hd5;
frames[2][3][24] = 8'hd5;
frames[2][3][25] = 8'hd5;
frames[2][3][26] = 8'hd5;
frames[2][3][27] = 8'hd1;
frames[2][3][28] = 8'hd1;
frames[2][3][29] = 8'hd1;
frames[2][3][30] = 8'hd1;
frames[2][3][31] = 8'hd1;
frames[2][3][32] = 8'hd1;
frames[2][3][33] = 8'hd5;
frames[2][3][34] = 8'hd1;
frames[2][3][35] = 8'hd1;
frames[2][3][36] = 8'hd1;
frames[2][3][37] = 8'hd1;
frames[2][3][38] = 8'hb1;
frames[2][3][39] = 8'had;
frames[2][4][0] = 8'had;
frames[2][4][1] = 8'hac;
frames[2][4][2] = 8'had;
frames[2][4][3] = 8'h8d;
frames[2][4][4] = 8'h8d;
frames[2][4][5] = 8'h8d;
frames[2][4][6] = 8'had;
frames[2][4][7] = 8'h89;
frames[2][4][8] = 8'had;
frames[2][4][9] = 8'hd1;
frames[2][4][10] = 8'hd1;
frames[2][4][11] = 8'hd1;
frames[2][4][12] = 8'hd5;
frames[2][4][13] = 8'hd5;
frames[2][4][14] = 8'hd5;
frames[2][4][15] = 8'hd5;
frames[2][4][16] = 8'hd1;
frames[2][4][17] = 8'hd1;
frames[2][4][18] = 8'hd1;
frames[2][4][19] = 8'hd1;
frames[2][4][20] = 8'hd1;
frames[2][4][21] = 8'hd1;
frames[2][4][22] = 8'hd5;
frames[2][4][23] = 8'hd5;
frames[2][4][24] = 8'hd5;
frames[2][4][25] = 8'hd5;
frames[2][4][26] = 8'hd5;
frames[2][4][27] = 8'hd5;
frames[2][4][28] = 8'hd1;
frames[2][4][29] = 8'hd1;
frames[2][4][30] = 8'hd1;
frames[2][4][31] = 8'hd1;
frames[2][4][32] = 8'hd1;
frames[2][4][33] = 8'hd5;
frames[2][4][34] = 8'hd5;
frames[2][4][35] = 8'hd1;
frames[2][4][36] = 8'hd1;
frames[2][4][37] = 8'hd1;
frames[2][4][38] = 8'hd1;
frames[2][4][39] = 8'had;
frames[2][5][0] = 8'hac;
frames[2][5][1] = 8'hac;
frames[2][5][2] = 8'had;
frames[2][5][3] = 8'had;
frames[2][5][4] = 8'h8d;
frames[2][5][5] = 8'h8d;
frames[2][5][6] = 8'had;
frames[2][5][7] = 8'h88;
frames[2][5][8] = 8'h68;
frames[2][5][9] = 8'hb1;
frames[2][5][10] = 8'hd1;
frames[2][5][11] = 8'hd1;
frames[2][5][12] = 8'hd1;
frames[2][5][13] = 8'hd1;
frames[2][5][14] = 8'hd1;
frames[2][5][15] = 8'hd1;
frames[2][5][16] = 8'hd1;
frames[2][5][17] = 8'hd1;
frames[2][5][18] = 8'hd1;
frames[2][5][19] = 8'hd1;
frames[2][5][20] = 8'hb1;
frames[2][5][21] = 8'hb1;
frames[2][5][22] = 8'hd1;
frames[2][5][23] = 8'hd1;
frames[2][5][24] = 8'hd5;
frames[2][5][25] = 8'hd5;
frames[2][5][26] = 8'hd5;
frames[2][5][27] = 8'hd5;
frames[2][5][28] = 8'hd1;
frames[2][5][29] = 8'hd1;
frames[2][5][30] = 8'hd1;
frames[2][5][31] = 8'hd1;
frames[2][5][32] = 8'hd1;
frames[2][5][33] = 8'hd5;
frames[2][5][34] = 8'hd5;
frames[2][5][35] = 8'hd1;
frames[2][5][36] = 8'hd1;
frames[2][5][37] = 8'hd1;
frames[2][5][38] = 8'hd1;
frames[2][5][39] = 8'had;
frames[2][6][0] = 8'hac;
frames[2][6][1] = 8'hac;
frames[2][6][2] = 8'hac;
frames[2][6][3] = 8'had;
frames[2][6][4] = 8'had;
frames[2][6][5] = 8'hac;
frames[2][6][6] = 8'h8d;
frames[2][6][7] = 8'had;
frames[2][6][8] = 8'h8d;
frames[2][6][9] = 8'hd1;
frames[2][6][10] = 8'hf6;
frames[2][6][11] = 8'hfa;
frames[2][6][12] = 8'hd6;
frames[2][6][13] = 8'hb1;
frames[2][6][14] = 8'hb1;
frames[2][6][15] = 8'hb1;
frames[2][6][16] = 8'hb1;
frames[2][6][17] = 8'h8d;
frames[2][6][18] = 8'h96;
frames[2][6][19] = 8'hb6;
frames[2][6][20] = 8'h96;
frames[2][6][21] = 8'h96;
frames[2][6][22] = 8'hb6;
frames[2][6][23] = 8'h92;
frames[2][6][24] = 8'h8d;
frames[2][6][25] = 8'h44;
frames[2][6][26] = 8'h8c;
frames[2][6][27] = 8'hd5;
frames[2][6][28] = 8'hd1;
frames[2][6][29] = 8'hd1;
frames[2][6][30] = 8'hd1;
frames[2][6][31] = 8'hd1;
frames[2][6][32] = 8'hd1;
frames[2][6][33] = 8'hd5;
frames[2][6][34] = 8'hd5;
frames[2][6][35] = 8'hd1;
frames[2][6][36] = 8'hd1;
frames[2][6][37] = 8'hd1;
frames[2][6][38] = 8'hd1;
frames[2][6][39] = 8'had;
frames[2][7][0] = 8'hac;
frames[2][7][1] = 8'hac;
frames[2][7][2] = 8'hac;
frames[2][7][3] = 8'hac;
frames[2][7][4] = 8'hac;
frames[2][7][5] = 8'hac;
frames[2][7][6] = 8'had;
frames[2][7][7] = 8'had;
frames[2][7][8] = 8'hd1;
frames[2][7][9] = 8'hfa;
frames[2][7][10] = 8'hfe;
frames[2][7][11] = 8'hfa;
frames[2][7][12] = 8'hfa;
frames[2][7][13] = 8'hb5;
frames[2][7][14] = 8'h8d;
frames[2][7][15] = 8'h8d;
frames[2][7][16] = 8'h6d;
frames[2][7][17] = 8'h91;
frames[2][7][18] = 8'hb6;
frames[2][7][19] = 8'h96;
frames[2][7][20] = 8'hda;
frames[2][7][21] = 8'hda;
frames[2][7][22] = 8'hda;
frames[2][7][23] = 8'hb6;
frames[2][7][24] = 8'h92;
frames[2][7][25] = 8'h24;
frames[2][7][26] = 8'h68;
frames[2][7][27] = 8'hd5;
frames[2][7][28] = 8'hd1;
frames[2][7][29] = 8'hd1;
frames[2][7][30] = 8'hd1;
frames[2][7][31] = 8'hd1;
frames[2][7][32] = 8'hd1;
frames[2][7][33] = 8'hd5;
frames[2][7][34] = 8'hd5;
frames[2][7][35] = 8'hd5;
frames[2][7][36] = 8'hd1;
frames[2][7][37] = 8'hd1;
frames[2][7][38] = 8'hd1;
frames[2][7][39] = 8'had;
frames[2][8][0] = 8'h8c;
frames[2][8][1] = 8'hac;
frames[2][8][2] = 8'hac;
frames[2][8][3] = 8'hac;
frames[2][8][4] = 8'hac;
frames[2][8][5] = 8'hac;
frames[2][8][6] = 8'h8d;
frames[2][8][7] = 8'hb1;
frames[2][8][8] = 8'hd6;
frames[2][8][9] = 8'hfa;
frames[2][8][10] = 8'hfa;
frames[2][8][11] = 8'hfa;
frames[2][8][12] = 8'hfa;
frames[2][8][13] = 8'hd6;
frames[2][8][14] = 8'h91;
frames[2][8][15] = 8'h8d;
frames[2][8][16] = 8'h91;
frames[2][8][17] = 8'hb6;
frames[2][8][18] = 8'hd6;
frames[2][8][19] = 8'hda;
frames[2][8][20] = 8'hfa;
frames[2][8][21] = 8'hfa;
frames[2][8][22] = 8'hfa;
frames[2][8][23] = 8'hfa;
frames[2][8][24] = 8'hb6;
frames[2][8][25] = 8'h91;
frames[2][8][26] = 8'h68;
frames[2][8][27] = 8'hd5;
frames[2][8][28] = 8'hd5;
frames[2][8][29] = 8'hd5;
frames[2][8][30] = 8'hd1;
frames[2][8][31] = 8'hd1;
frames[2][8][32] = 8'hd1;
frames[2][8][33] = 8'hd5;
frames[2][8][34] = 8'hd5;
frames[2][8][35] = 8'hd5;
frames[2][8][36] = 8'hd1;
frames[2][8][37] = 8'hd1;
frames[2][8][38] = 8'hd1;
frames[2][8][39] = 8'had;
frames[2][9][0] = 8'h8c;
frames[2][9][1] = 8'hac;
frames[2][9][2] = 8'hac;
frames[2][9][3] = 8'had;
frames[2][9][4] = 8'hac;
frames[2][9][5] = 8'hac;
frames[2][9][6] = 8'h8d;
frames[2][9][7] = 8'h8d;
frames[2][9][8] = 8'hb1;
frames[2][9][9] = 8'hfa;
frames[2][9][10] = 8'hfa;
frames[2][9][11] = 8'hfa;
frames[2][9][12] = 8'hfa;
frames[2][9][13] = 8'hd6;
frames[2][9][14] = 8'h91;
frames[2][9][15] = 8'h91;
frames[2][9][16] = 8'hb6;
frames[2][9][17] = 8'hda;
frames[2][9][18] = 8'hfa;
frames[2][9][19] = 8'hfa;
frames[2][9][20] = 8'hfa;
frames[2][9][21] = 8'hfa;
frames[2][9][22] = 8'hfa;
frames[2][9][23] = 8'hfa;
frames[2][9][24] = 8'hfb;
frames[2][9][25] = 8'hb6;
frames[2][9][26] = 8'hb1;
frames[2][9][27] = 8'hb5;
frames[2][9][28] = 8'hd5;
frames[2][9][29] = 8'hd1;
frames[2][9][30] = 8'hd1;
frames[2][9][31] = 8'hd1;
frames[2][9][32] = 8'hd1;
frames[2][9][33] = 8'hd5;
frames[2][9][34] = 8'hd5;
frames[2][9][35] = 8'hd5;
frames[2][9][36] = 8'hd1;
frames[2][9][37] = 8'hd1;
frames[2][9][38] = 8'hd1;
frames[2][9][39] = 8'hb1;
frames[2][10][0] = 8'hac;
frames[2][10][1] = 8'hac;
frames[2][10][2] = 8'hac;
frames[2][10][3] = 8'hac;
frames[2][10][4] = 8'hac;
frames[2][10][5] = 8'hac;
frames[2][10][6] = 8'h8c;
frames[2][10][7] = 8'h8c;
frames[2][10][8] = 8'hb5;
frames[2][10][9] = 8'hfa;
frames[2][10][10] = 8'hfa;
frames[2][10][11] = 8'hfa;
frames[2][10][12] = 8'hfa;
frames[2][10][13] = 8'hd6;
frames[2][10][14] = 8'h91;
frames[2][10][15] = 8'hb2;
frames[2][10][16] = 8'hfa;
frames[2][10][17] = 8'hfb;
frames[2][10][18] = 8'hfa;
frames[2][10][19] = 8'hfa;
frames[2][10][20] = 8'hfa;
frames[2][10][21] = 8'hfa;
frames[2][10][22] = 8'hfa;
frames[2][10][23] = 8'hfa;
frames[2][10][24] = 8'hfa;
frames[2][10][25] = 8'hfa;
frames[2][10][26] = 8'hd6;
frames[2][10][27] = 8'hb5;
frames[2][10][28] = 8'hd5;
frames[2][10][29] = 8'hd1;
frames[2][10][30] = 8'hd1;
frames[2][10][31] = 8'hd1;
frames[2][10][32] = 8'hd1;
frames[2][10][33] = 8'hd1;
frames[2][10][34] = 8'hd5;
frames[2][10][35] = 8'hd5;
frames[2][10][36] = 8'hd1;
frames[2][10][37] = 8'hd1;
frames[2][10][38] = 8'hd1;
frames[2][10][39] = 8'hb1;
frames[2][11][0] = 8'hac;
frames[2][11][1] = 8'hac;
frames[2][11][2] = 8'hac;
frames[2][11][3] = 8'hac;
frames[2][11][4] = 8'hac;
frames[2][11][5] = 8'hac;
frames[2][11][6] = 8'h8c;
frames[2][11][7] = 8'h8c;
frames[2][11][8] = 8'hd5;
frames[2][11][9] = 8'hd6;
frames[2][11][10] = 8'hfa;
frames[2][11][11] = 8'hfa;
frames[2][11][12] = 8'hda;
frames[2][11][13] = 8'hb5;
frames[2][11][14] = 8'hb1;
frames[2][11][15] = 8'hd6;
frames[2][11][16] = 8'hfa;
frames[2][11][17] = 8'hfb;
frames[2][11][18] = 8'hfb;
frames[2][11][19] = 8'hfa;
frames[2][11][20] = 8'hfa;
frames[2][11][21] = 8'hfa;
frames[2][11][22] = 8'hfa;
frames[2][11][23] = 8'hfa;
frames[2][11][24] = 8'hfa;
frames[2][11][25] = 8'hfa;
frames[2][11][26] = 8'hda;
frames[2][11][27] = 8'hb5;
frames[2][11][28] = 8'hd1;
frames[2][11][29] = 8'hd1;
frames[2][11][30] = 8'hd1;
frames[2][11][31] = 8'hd1;
frames[2][11][32] = 8'hd1;
frames[2][11][33] = 8'hd1;
frames[2][11][34] = 8'hd5;
frames[2][11][35] = 8'hd5;
frames[2][11][36] = 8'hd1;
frames[2][11][37] = 8'hd1;
frames[2][11][38] = 8'hd1;
frames[2][11][39] = 8'hb1;
frames[2][12][0] = 8'h8c;
frames[2][12][1] = 8'hac;
frames[2][12][2] = 8'hac;
frames[2][12][3] = 8'hac;
frames[2][12][4] = 8'hac;
frames[2][12][5] = 8'hac;
frames[2][12][6] = 8'h8c;
frames[2][12][7] = 8'h88;
frames[2][12][8] = 8'hb1;
frames[2][12][9] = 8'hd6;
frames[2][12][10] = 8'hfa;
frames[2][12][11] = 8'hfa;
frames[2][12][12] = 8'hda;
frames[2][12][13] = 8'h91;
frames[2][12][14] = 8'hb1;
frames[2][12][15] = 8'hda;
frames[2][12][16] = 8'hfb;
frames[2][12][17] = 8'hfb;
frames[2][12][18] = 8'hfa;
frames[2][12][19] = 8'hfa;
frames[2][12][20] = 8'hfa;
frames[2][12][21] = 8'hfa;
frames[2][12][22] = 8'hfa;
frames[2][12][23] = 8'hfa;
frames[2][12][24] = 8'hfa;
frames[2][12][25] = 8'hfa;
frames[2][12][26] = 8'hfa;
frames[2][12][27] = 8'hb6;
frames[2][12][28] = 8'hd1;
frames[2][12][29] = 8'hd5;
frames[2][12][30] = 8'hd1;
frames[2][12][31] = 8'hd1;
frames[2][12][32] = 8'hd1;
frames[2][12][33] = 8'hd1;
frames[2][12][34] = 8'hd5;
frames[2][12][35] = 8'hd5;
frames[2][12][36] = 8'hd1;
frames[2][12][37] = 8'hd1;
frames[2][12][38] = 8'hd1;
frames[2][12][39] = 8'hb1;
frames[2][13][0] = 8'h8c;
frames[2][13][1] = 8'h8c;
frames[2][13][2] = 8'hac;
frames[2][13][3] = 8'hac;
frames[2][13][4] = 8'hac;
frames[2][13][5] = 8'hac;
frames[2][13][6] = 8'h8c;
frames[2][13][7] = 8'h8c;
frames[2][13][8] = 8'h91;
frames[2][13][9] = 8'hb5;
frames[2][13][10] = 8'hda;
frames[2][13][11] = 8'hfa;
frames[2][13][12] = 8'hb1;
frames[2][13][13] = 8'h8d;
frames[2][13][14] = 8'h91;
frames[2][13][15] = 8'hda;
frames[2][13][16] = 8'hfb;
frames[2][13][17] = 8'hfb;
frames[2][13][18] = 8'hfa;
frames[2][13][19] = 8'hfa;
frames[2][13][20] = 8'hfa;
frames[2][13][21] = 8'hfa;
frames[2][13][22] = 8'hfa;
frames[2][13][23] = 8'hfa;
frames[2][13][24] = 8'hfa;
frames[2][13][25] = 8'hfa;
frames[2][13][26] = 8'hfa;
frames[2][13][27] = 8'hd6;
frames[2][13][28] = 8'hd1;
frames[2][13][29] = 8'hd5;
frames[2][13][30] = 8'hd1;
frames[2][13][31] = 8'hd1;
frames[2][13][32] = 8'hd1;
frames[2][13][33] = 8'hd1;
frames[2][13][34] = 8'hd5;
frames[2][13][35] = 8'hd5;
frames[2][13][36] = 8'hd1;
frames[2][13][37] = 8'hd1;
frames[2][13][38] = 8'hb1;
frames[2][13][39] = 8'hb1;
frames[2][14][0] = 8'h8c;
frames[2][14][1] = 8'hac;
frames[2][14][2] = 8'hac;
frames[2][14][3] = 8'hac;
frames[2][14][4] = 8'hac;
frames[2][14][5] = 8'hac;
frames[2][14][6] = 8'h8c;
frames[2][14][7] = 8'h68;
frames[2][14][8] = 8'h8d;
frames[2][14][9] = 8'h91;
frames[2][14][10] = 8'hb1;
frames[2][14][11] = 8'h8d;
frames[2][14][12] = 8'h8d;
frames[2][14][13] = 8'h8d;
frames[2][14][14] = 8'h8d;
frames[2][14][15] = 8'hd6;
frames[2][14][16] = 8'hff;
frames[2][14][17] = 8'hff;
frames[2][14][18] = 8'hfb;
frames[2][14][19] = 8'hfa;
frames[2][14][20] = 8'hfa;
frames[2][14][21] = 8'hfa;
frames[2][14][22] = 8'hfa;
frames[2][14][23] = 8'hfa;
frames[2][14][24] = 8'hfb;
frames[2][14][25] = 8'hfb;
frames[2][14][26] = 8'hfa;
frames[2][14][27] = 8'hd6;
frames[2][14][28] = 8'hd1;
frames[2][14][29] = 8'hd5;
frames[2][14][30] = 8'hd1;
frames[2][14][31] = 8'hd1;
frames[2][14][32] = 8'hd1;
frames[2][14][33] = 8'hd1;
frames[2][14][34] = 8'hd1;
frames[2][14][35] = 8'hd5;
frames[2][14][36] = 8'hd1;
frames[2][14][37] = 8'hd1;
frames[2][14][38] = 8'hb1;
frames[2][14][39] = 8'hb1;
frames[2][15][0] = 8'h8c;
frames[2][15][1] = 8'hac;
frames[2][15][2] = 8'hac;
frames[2][15][3] = 8'hac;
frames[2][15][4] = 8'hac;
frames[2][15][5] = 8'hac;
frames[2][15][6] = 8'h88;
frames[2][15][7] = 8'h68;
frames[2][15][8] = 8'h89;
frames[2][15][9] = 8'h68;
frames[2][15][10] = 8'h69;
frames[2][15][11] = 8'h8d;
frames[2][15][12] = 8'h8d;
frames[2][15][13] = 8'h8d;
frames[2][15][14] = 8'h8d;
frames[2][15][15] = 8'hb6;
frames[2][15][16] = 8'hfb;
frames[2][15][17] = 8'hff;
frames[2][15][18] = 8'hfb;
frames[2][15][19] = 8'hfb;
frames[2][15][20] = 8'hfa;
frames[2][15][21] = 8'hfa;
frames[2][15][22] = 8'hfa;
frames[2][15][23] = 8'hfa;
frames[2][15][24] = 8'hfb;
frames[2][15][25] = 8'hfb;
frames[2][15][26] = 8'hda;
frames[2][15][27] = 8'hb6;
frames[2][15][28] = 8'hd1;
frames[2][15][29] = 8'hd1;
frames[2][15][30] = 8'hd1;
frames[2][15][31] = 8'hd1;
frames[2][15][32] = 8'hd1;
frames[2][15][33] = 8'hd1;
frames[2][15][34] = 8'hd1;
frames[2][15][35] = 8'hd1;
frames[2][15][36] = 8'hd1;
frames[2][15][37] = 8'hd1;
frames[2][15][38] = 8'hb1;
frames[2][15][39] = 8'hb1;
frames[2][16][0] = 8'h8c;
frames[2][16][1] = 8'h8c;
frames[2][16][2] = 8'h8c;
frames[2][16][3] = 8'h8c;
frames[2][16][4] = 8'h8c;
frames[2][16][5] = 8'h8c;
frames[2][16][6] = 8'h88;
frames[2][16][7] = 8'h88;
frames[2][16][8] = 8'h88;
frames[2][16][9] = 8'h40;
frames[2][16][10] = 8'h64;
frames[2][16][11] = 8'h89;
frames[2][16][12] = 8'h8d;
frames[2][16][13] = 8'h8d;
frames[2][16][14] = 8'h8d;
frames[2][16][15] = 8'h91;
frames[2][16][16] = 8'hfa;
frames[2][16][17] = 8'hfb;
frames[2][16][18] = 8'hfa;
frames[2][16][19] = 8'hfa;
frames[2][16][20] = 8'hfa;
frames[2][16][21] = 8'hfa;
frames[2][16][22] = 8'hfa;
frames[2][16][23] = 8'hfb;
frames[2][16][24] = 8'hfb;
frames[2][16][25] = 8'hfb;
frames[2][16][26] = 8'hd6;
frames[2][16][27] = 8'hb1;
frames[2][16][28] = 8'hd1;
frames[2][16][29] = 8'hd1;
frames[2][16][30] = 8'hd1;
frames[2][16][31] = 8'hd1;
frames[2][16][32] = 8'hd1;
frames[2][16][33] = 8'hd1;
frames[2][16][34] = 8'hd1;
frames[2][16][35] = 8'hd1;
frames[2][16][36] = 8'hd1;
frames[2][16][37] = 8'hb1;
frames[2][16][38] = 8'hb1;
frames[2][16][39] = 8'hb1;
frames[2][17][0] = 8'h8c;
frames[2][17][1] = 8'h8c;
frames[2][17][2] = 8'h8c;
frames[2][17][3] = 8'h8c;
frames[2][17][4] = 8'h8c;
frames[2][17][5] = 8'h8c;
frames[2][17][6] = 8'h88;
frames[2][17][7] = 8'h68;
frames[2][17][8] = 8'h60;
frames[2][17][9] = 8'h40;
frames[2][17][10] = 8'h40;
frames[2][17][11] = 8'h64;
frames[2][17][12] = 8'h8d;
frames[2][17][13] = 8'h8d;
frames[2][17][14] = 8'h8d;
frames[2][17][15] = 8'h8d;
frames[2][17][16] = 8'hd6;
frames[2][17][17] = 8'hfb;
frames[2][17][18] = 8'hfa;
frames[2][17][19] = 8'hfa;
frames[2][17][20] = 8'hfa;
frames[2][17][21] = 8'hfa;
frames[2][17][22] = 8'hfb;
frames[2][17][23] = 8'hfa;
frames[2][17][24] = 8'hfb;
frames[2][17][25] = 8'hfb;
frames[2][17][26] = 8'hb1;
frames[2][17][27] = 8'h6d;
frames[2][17][28] = 8'hd1;
frames[2][17][29] = 8'hd1;
frames[2][17][30] = 8'hd1;
frames[2][17][31] = 8'hd1;
frames[2][17][32] = 8'hd1;
frames[2][17][33] = 8'hd1;
frames[2][17][34] = 8'hd1;
frames[2][17][35] = 8'hd1;
frames[2][17][36] = 8'hd1;
frames[2][17][37] = 8'hb1;
frames[2][17][38] = 8'hb1;
frames[2][17][39] = 8'hb1;
frames[2][18][0] = 8'h8c;
frames[2][18][1] = 8'h8c;
frames[2][18][2] = 8'hac;
frames[2][18][3] = 8'hac;
frames[2][18][4] = 8'hac;
frames[2][18][5] = 8'h8c;
frames[2][18][6] = 8'h68;
frames[2][18][7] = 8'h64;
frames[2][18][8] = 8'h40;
frames[2][18][9] = 8'h40;
frames[2][18][10] = 8'h40;
frames[2][18][11] = 8'h64;
frames[2][18][12] = 8'h69;
frames[2][18][13] = 8'h8d;
frames[2][18][14] = 8'h8d;
frames[2][18][15] = 8'h8d;
frames[2][18][16] = 8'h91;
frames[2][18][17] = 8'hda;
frames[2][18][18] = 8'hfa;
frames[2][18][19] = 8'hfa;
frames[2][18][20] = 8'hfa;
frames[2][18][21] = 8'hfa;
frames[2][18][22] = 8'hfa;
frames[2][18][23] = 8'hfa;
frames[2][18][24] = 8'hfb;
frames[2][18][25] = 8'hda;
frames[2][18][26] = 8'h8d;
frames[2][18][27] = 8'h6d;
frames[2][18][28] = 8'hd1;
frames[2][18][29] = 8'hd1;
frames[2][18][30] = 8'hd1;
frames[2][18][31] = 8'hd1;
frames[2][18][32] = 8'hd1;
frames[2][18][33] = 8'hd1;
frames[2][18][34] = 8'hd1;
frames[2][18][35] = 8'hd1;
frames[2][18][36] = 8'hd1;
frames[2][18][37] = 8'hb1;
frames[2][18][38] = 8'hb1;
frames[2][18][39] = 8'hb1;
frames[2][19][0] = 8'h8c;
frames[2][19][1] = 8'h8c;
frames[2][19][2] = 8'hac;
frames[2][19][3] = 8'hac;
frames[2][19][4] = 8'hac;
frames[2][19][5] = 8'h8c;
frames[2][19][6] = 8'h68;
frames[2][19][7] = 8'h64;
frames[2][19][8] = 8'h40;
frames[2][19][9] = 8'h40;
frames[2][19][10] = 8'h40;
frames[2][19][11] = 8'h64;
frames[2][19][12] = 8'h68;
frames[2][19][13] = 8'h6d;
frames[2][19][14] = 8'h89;
frames[2][19][15] = 8'h69;
frames[2][19][16] = 8'h69;
frames[2][19][17] = 8'hb2;
frames[2][19][18] = 8'hda;
frames[2][19][19] = 8'hda;
frames[2][19][20] = 8'hda;
frames[2][19][21] = 8'hda;
frames[2][19][22] = 8'hda;
frames[2][19][23] = 8'hfa;
frames[2][19][24] = 8'hda;
frames[2][19][25] = 8'hb6;
frames[2][19][26] = 8'h6d;
frames[2][19][27] = 8'h6d;
frames[2][19][28] = 8'hd1;
frames[2][19][29] = 8'hd1;
frames[2][19][30] = 8'hd1;
frames[2][19][31] = 8'hd1;
frames[2][19][32] = 8'hd1;
frames[2][19][33] = 8'hd1;
frames[2][19][34] = 8'hd1;
frames[2][19][35] = 8'hd1;
frames[2][19][36] = 8'hd1;
frames[2][19][37] = 8'hb1;
frames[2][19][38] = 8'hb1;
frames[2][19][39] = 8'hb1;
frames[2][20][0] = 8'h8c;
frames[2][20][1] = 8'h8c;
frames[2][20][2] = 8'h8c;
frames[2][20][3] = 8'h8c;
frames[2][20][4] = 8'h8c;
frames[2][20][5] = 8'h8c;
frames[2][20][6] = 8'h68;
frames[2][20][7] = 8'h88;
frames[2][20][8] = 8'h68;
frames[2][20][9] = 8'h64;
frames[2][20][10] = 8'h68;
frames[2][20][11] = 8'h68;
frames[2][20][12] = 8'h68;
frames[2][20][13] = 8'h8d;
frames[2][20][14] = 8'h88;
frames[2][20][15] = 8'h88;
frames[2][20][16] = 8'h88;
frames[2][20][17] = 8'h88;
frames[2][20][18] = 8'hb6;
frames[2][20][19] = 8'hba;
frames[2][20][20] = 8'hb6;
frames[2][20][21] = 8'hb6;
frames[2][20][22] = 8'hba;
frames[2][20][23] = 8'hda;
frames[2][20][24] = 8'hb6;
frames[2][20][25] = 8'h91;
frames[2][20][26] = 8'h6d;
frames[2][20][27] = 8'h69;
frames[2][20][28] = 8'hd1;
frames[2][20][29] = 8'hd1;
frames[2][20][30] = 8'hd1;
frames[2][20][31] = 8'hd1;
frames[2][20][32] = 8'hd1;
frames[2][20][33] = 8'hd1;
frames[2][20][34] = 8'hd1;
frames[2][20][35] = 8'hd1;
frames[2][20][36] = 8'hb1;
frames[2][20][37] = 8'hb1;
frames[2][20][38] = 8'hb1;
frames[2][20][39] = 8'hb1;
frames[2][21][0] = 8'h88;
frames[2][21][1] = 8'h88;
frames[2][21][2] = 8'h88;
frames[2][21][3] = 8'h88;
frames[2][21][4] = 8'h88;
frames[2][21][5] = 8'h88;
frames[2][21][6] = 8'h68;
frames[2][21][7] = 8'h8d;
frames[2][21][8] = 8'h8d;
frames[2][21][9] = 8'h69;
frames[2][21][10] = 8'h69;
frames[2][21][11] = 8'h69;
frames[2][21][12] = 8'h69;
frames[2][21][13] = 8'h8d;
frames[2][21][14] = 8'h84;
frames[2][21][15] = 8'h84;
frames[2][21][16] = 8'h84;
frames[2][21][17] = 8'h84;
frames[2][21][18] = 8'h8d;
frames[2][21][19] = 8'h92;
frames[2][21][20] = 8'hb6;
frames[2][21][21] = 8'hb6;
frames[2][21][22] = 8'hb6;
frames[2][21][23] = 8'hb2;
frames[2][21][24] = 8'h91;
frames[2][21][25] = 8'h91;
frames[2][21][26] = 8'h6d;
frames[2][21][27] = 8'h68;
frames[2][21][28] = 8'hd1;
frames[2][21][29] = 8'hd1;
frames[2][21][30] = 8'hd1;
frames[2][21][31] = 8'hd1;
frames[2][21][32] = 8'hd1;
frames[2][21][33] = 8'hd1;
frames[2][21][34] = 8'hb1;
frames[2][21][35] = 8'hd1;
frames[2][21][36] = 8'hb1;
frames[2][21][37] = 8'hb1;
frames[2][21][38] = 8'hb1;
frames[2][21][39] = 8'hb1;
frames[2][22][0] = 8'h88;
frames[2][22][1] = 8'h88;
frames[2][22][2] = 8'h88;
frames[2][22][3] = 8'h68;
frames[2][22][4] = 8'h68;
frames[2][22][5] = 8'h68;
frames[2][22][6] = 8'h64;
frames[2][22][7] = 8'h8d;
frames[2][22][8] = 8'h69;
frames[2][22][9] = 8'h6d;
frames[2][22][10] = 8'h6d;
frames[2][22][11] = 8'h6d;
frames[2][22][12] = 8'h8d;
frames[2][22][13] = 8'h8d;
frames[2][22][14] = 8'h84;
frames[2][22][15] = 8'h84;
frames[2][22][16] = 8'ha8;
frames[2][22][17] = 8'ha8;
frames[2][22][18] = 8'h91;
frames[2][22][19] = 8'h8d;
frames[2][22][20] = 8'h8d;
frames[2][22][21] = 8'h8d;
frames[2][22][22] = 8'h8d;
frames[2][22][23] = 8'h91;
frames[2][22][24] = 8'h91;
frames[2][22][25] = 8'h91;
frames[2][22][26] = 8'h68;
frames[2][22][27] = 8'h44;
frames[2][22][28] = 8'hd1;
frames[2][22][29] = 8'hd1;
frames[2][22][30] = 8'hd1;
frames[2][22][31] = 8'hd1;
frames[2][22][32] = 8'hd1;
frames[2][22][33] = 8'hd1;
frames[2][22][34] = 8'hb1;
frames[2][22][35] = 8'hd1;
frames[2][22][36] = 8'hb1;
frames[2][22][37] = 8'hb1;
frames[2][22][38] = 8'hb1;
frames[2][22][39] = 8'hb1;
frames[2][23][0] = 8'h88;
frames[2][23][1] = 8'h88;
frames[2][23][2] = 8'h68;
frames[2][23][3] = 8'h68;
frames[2][23][4] = 8'h68;
frames[2][23][5] = 8'h88;
frames[2][23][6] = 8'h88;
frames[2][23][7] = 8'h88;
frames[2][23][8] = 8'h44;
frames[2][23][9] = 8'h69;
frames[2][23][10] = 8'h89;
frames[2][23][11] = 8'h89;
frames[2][23][12] = 8'h6d;
frames[2][23][13] = 8'h8d;
frames[2][23][14] = 8'h88;
frames[2][23][15] = 8'h64;
frames[2][23][16] = 8'h64;
frames[2][23][17] = 8'h88;
frames[2][23][18] = 8'h8d;
frames[2][23][19] = 8'h6d;
frames[2][23][20] = 8'h69;
frames[2][23][21] = 8'h69;
frames[2][23][22] = 8'h69;
frames[2][23][23] = 8'h69;
frames[2][23][24] = 8'h68;
frames[2][23][25] = 8'h48;
frames[2][23][26] = 8'h24;
frames[2][23][27] = 8'h69;
frames[2][23][28] = 8'hd5;
frames[2][23][29] = 8'hd1;
frames[2][23][30] = 8'hd1;
frames[2][23][31] = 8'hd1;
frames[2][23][32] = 8'hd1;
frames[2][23][33] = 8'hb1;
frames[2][23][34] = 8'hb1;
frames[2][23][35] = 8'hd1;
frames[2][23][36] = 8'hb1;
frames[2][23][37] = 8'hb1;
frames[2][23][38] = 8'hb1;
frames[2][23][39] = 8'hb1;
frames[2][24][0] = 8'h68;
frames[2][24][1] = 8'h68;
frames[2][24][2] = 8'h88;
frames[2][24][3] = 8'h8d;
frames[2][24][4] = 8'hd1;
frames[2][24][5] = 8'hd1;
frames[2][24][6] = 8'hd1;
frames[2][24][7] = 8'had;
frames[2][24][8] = 8'had;
frames[2][24][9] = 8'h89;
frames[2][24][10] = 8'h44;
frames[2][24][11] = 8'h44;
frames[2][24][12] = 8'h44;
frames[2][24][13] = 8'h8d;
frames[2][24][14] = 8'h8d;
frames[2][24][15] = 8'h44;
frames[2][24][16] = 8'h68;
frames[2][24][17] = 8'h68;
frames[2][24][18] = 8'h8d;
frames[2][24][19] = 8'h8d;
frames[2][24][20] = 8'h8d;
frames[2][24][21] = 8'h8d;
frames[2][24][22] = 8'h8d;
frames[2][24][23] = 8'h8d;
frames[2][24][24] = 8'h91;
frames[2][24][25] = 8'hb1;
frames[2][24][26] = 8'hb1;
frames[2][24][27] = 8'hb5;
frames[2][24][28] = 8'hd1;
frames[2][24][29] = 8'hd1;
frames[2][24][30] = 8'hd1;
frames[2][24][31] = 8'hd1;
frames[2][24][32] = 8'hb1;
frames[2][24][33] = 8'hb1;
frames[2][24][34] = 8'hb1;
frames[2][24][35] = 8'hd1;
frames[2][24][36] = 8'hb1;
frames[2][24][37] = 8'hb1;
frames[2][24][38] = 8'hb1;
frames[2][24][39] = 8'hb1;
frames[2][25][0] = 8'had;
frames[2][25][1] = 8'hd1;
frames[2][25][2] = 8'hd1;
frames[2][25][3] = 8'hd1;
frames[2][25][4] = 8'hd1;
frames[2][25][5] = 8'hb1;
frames[2][25][6] = 8'hd1;
frames[2][25][7] = 8'h88;
frames[2][25][8] = 8'h44;
frames[2][25][9] = 8'h89;
frames[2][25][10] = 8'h8d;
frames[2][25][11] = 8'h8d;
frames[2][25][12] = 8'h8d;
frames[2][25][13] = 8'hb1;
frames[2][25][14] = 8'hb1;
frames[2][25][15] = 8'hb1;
frames[2][25][16] = 8'hb1;
frames[2][25][17] = 8'hb1;
frames[2][25][18] = 8'hb1;
frames[2][25][19] = 8'hd1;
frames[2][25][20] = 8'hd5;
frames[2][25][21] = 8'hd1;
frames[2][25][22] = 8'hd1;
frames[2][25][23] = 8'hd5;
frames[2][25][24] = 8'hd1;
frames[2][25][25] = 8'hd1;
frames[2][25][26] = 8'hd1;
frames[2][25][27] = 8'hd1;
frames[2][25][28] = 8'hd1;
frames[2][25][29] = 8'hd1;
frames[2][25][30] = 8'hd1;
frames[2][25][31] = 8'hd1;
frames[2][25][32] = 8'hb1;
frames[2][25][33] = 8'hb1;
frames[2][25][34] = 8'hb1;
frames[2][25][35] = 8'hb1;
frames[2][25][36] = 8'hb1;
frames[2][25][37] = 8'hb1;
frames[2][25][38] = 8'hb1;
frames[2][25][39] = 8'hb1;
frames[2][26][0] = 8'had;
frames[2][26][1] = 8'had;
frames[2][26][2] = 8'had;
frames[2][26][3] = 8'had;
frames[2][26][4] = 8'had;
frames[2][26][5] = 8'had;
frames[2][26][6] = 8'hd1;
frames[2][26][7] = 8'had;
frames[2][26][8] = 8'h88;
frames[2][26][9] = 8'had;
frames[2][26][10] = 8'had;
frames[2][26][11] = 8'hb1;
frames[2][26][12] = 8'hb1;
frames[2][26][13] = 8'hb1;
frames[2][26][14] = 8'hb1;
frames[2][26][15] = 8'hb1;
frames[2][26][16] = 8'had;
frames[2][26][17] = 8'had;
frames[2][26][18] = 8'hb1;
frames[2][26][19] = 8'hb1;
frames[2][26][20] = 8'hd1;
frames[2][26][21] = 8'hd1;
frames[2][26][22] = 8'hd1;
frames[2][26][23] = 8'hd1;
frames[2][26][24] = 8'hd1;
frames[2][26][25] = 8'hd1;
frames[2][26][26] = 8'hd1;
frames[2][26][27] = 8'hd1;
frames[2][26][28] = 8'hd1;
frames[2][26][29] = 8'hb1;
frames[2][26][30] = 8'hb1;
frames[2][26][31] = 8'hb1;
frames[2][26][32] = 8'hb1;
frames[2][26][33] = 8'hb1;
frames[2][26][34] = 8'hb1;
frames[2][26][35] = 8'hb1;
frames[2][26][36] = 8'hb1;
frames[2][26][37] = 8'hb1;
frames[2][26][38] = 8'hb1;
frames[2][26][39] = 8'hb1;
frames[2][27][0] = 8'h88;
frames[2][27][1] = 8'h88;
frames[2][27][2] = 8'h88;
frames[2][27][3] = 8'h88;
frames[2][27][4] = 8'h88;
frames[2][27][5] = 8'h8d;
frames[2][27][6] = 8'had;
frames[2][27][7] = 8'hb1;
frames[2][27][8] = 8'had;
frames[2][27][9] = 8'had;
frames[2][27][10] = 8'had;
frames[2][27][11] = 8'hb1;
frames[2][27][12] = 8'hb1;
frames[2][27][13] = 8'hb1;
frames[2][27][14] = 8'hb1;
frames[2][27][15] = 8'hb1;
frames[2][27][16] = 8'hac;
frames[2][27][17] = 8'hac;
frames[2][27][18] = 8'hac;
frames[2][27][19] = 8'hb1;
frames[2][27][20] = 8'hb1;
frames[2][27][21] = 8'hd1;
frames[2][27][22] = 8'hd1;
frames[2][27][23] = 8'hd1;
frames[2][27][24] = 8'hd1;
frames[2][27][25] = 8'hd1;
frames[2][27][26] = 8'hd1;
frames[2][27][27] = 8'hb1;
frames[2][27][28] = 8'hb1;
frames[2][27][29] = 8'hb1;
frames[2][27][30] = 8'hb1;
frames[2][27][31] = 8'hb1;
frames[2][27][32] = 8'hb1;
frames[2][27][33] = 8'hb1;
frames[2][27][34] = 8'hb1;
frames[2][27][35] = 8'hb1;
frames[2][27][36] = 8'hb1;
frames[2][27][37] = 8'hb1;
frames[2][27][38] = 8'hb1;
frames[2][27][39] = 8'hb1;
frames[2][28][0] = 8'h88;
frames[2][28][1] = 8'h88;
frames[2][28][2] = 8'h68;
frames[2][28][3] = 8'h68;
frames[2][28][4] = 8'h88;
frames[2][28][5] = 8'h88;
frames[2][28][6] = 8'h88;
frames[2][28][7] = 8'had;
frames[2][28][8] = 8'had;
frames[2][28][9] = 8'had;
frames[2][28][10] = 8'hb1;
frames[2][28][11] = 8'hb1;
frames[2][28][12] = 8'hb1;
frames[2][28][13] = 8'hb1;
frames[2][28][14] = 8'hb1;
frames[2][28][15] = 8'hb1;
frames[2][28][16] = 8'hac;
frames[2][28][17] = 8'h8c;
frames[2][28][18] = 8'h8c;
frames[2][28][19] = 8'hac;
frames[2][28][20] = 8'hac;
frames[2][28][21] = 8'hb1;
frames[2][28][22] = 8'hd1;
frames[2][28][23] = 8'hd1;
frames[2][28][24] = 8'hd1;
frames[2][28][25] = 8'hd1;
frames[2][28][26] = 8'hb1;
frames[2][28][27] = 8'hb1;
frames[2][28][28] = 8'hb1;
frames[2][28][29] = 8'hb1;
frames[2][28][30] = 8'hb1;
frames[2][28][31] = 8'hb1;
frames[2][28][32] = 8'hb1;
frames[2][28][33] = 8'hb1;
frames[2][28][34] = 8'hb1;
frames[2][28][35] = 8'hb1;
frames[2][28][36] = 8'hb1;
frames[2][28][37] = 8'hb1;
frames[2][28][38] = 8'hb1;
frames[2][28][39] = 8'hb1;
frames[2][29][0] = 8'h68;
frames[2][29][1] = 8'h68;
frames[2][29][2] = 8'h68;
frames[2][29][3] = 8'h68;
frames[2][29][4] = 8'h88;
frames[2][29][5] = 8'h88;
frames[2][29][6] = 8'h88;
frames[2][29][7] = 8'h8d;
frames[2][29][8] = 8'had;
frames[2][29][9] = 8'had;
frames[2][29][10] = 8'hb1;
frames[2][29][11] = 8'hb1;
frames[2][29][12] = 8'hb1;
frames[2][29][13] = 8'hb1;
frames[2][29][14] = 8'hb1;
frames[2][29][15] = 8'hb1;
frames[2][29][16] = 8'hac;
frames[2][29][17] = 8'h8c;
frames[2][29][18] = 8'h8c;
frames[2][29][19] = 8'h8c;
frames[2][29][20] = 8'h8c;
frames[2][29][21] = 8'hac;
frames[2][29][22] = 8'hb1;
frames[2][29][23] = 8'hd1;
frames[2][29][24] = 8'hd1;
frames[2][29][25] = 8'hb1;
frames[2][29][26] = 8'hb1;
frames[2][29][27] = 8'hb1;
frames[2][29][28] = 8'hb1;
frames[2][29][29] = 8'hb1;
frames[2][29][30] = 8'hb1;
frames[2][29][31] = 8'hb1;
frames[2][29][32] = 8'hb1;
frames[2][29][33] = 8'hb1;
frames[2][29][34] = 8'hb1;
frames[2][29][35] = 8'hb1;
frames[2][29][36] = 8'hb1;
frames[2][29][37] = 8'hb1;
frames[2][29][38] = 8'hb1;
frames[2][29][39] = 8'hb1;
frames[3][0][0] = 8'hd1;
frames[3][0][1] = 8'hb1;
frames[3][0][2] = 8'hb1;
frames[3][0][3] = 8'hd1;
frames[3][0][4] = 8'hd1;
frames[3][0][5] = 8'hd1;
frames[3][0][6] = 8'hd1;
frames[3][0][7] = 8'hd5;
frames[3][0][8] = 8'hd5;
frames[3][0][9] = 8'hd1;
frames[3][0][10] = 8'hd1;
frames[3][0][11] = 8'hd5;
frames[3][0][12] = 8'hd5;
frames[3][0][13] = 8'hd5;
frames[3][0][14] = 8'hd5;
frames[3][0][15] = 8'hd5;
frames[3][0][16] = 8'hd5;
frames[3][0][17] = 8'hd1;
frames[3][0][18] = 8'hd5;
frames[3][0][19] = 8'hd1;
frames[3][0][20] = 8'hd1;
frames[3][0][21] = 8'hd1;
frames[3][0][22] = 8'hd5;
frames[3][0][23] = 8'hd5;
frames[3][0][24] = 8'hd5;
frames[3][0][25] = 8'hd5;
frames[3][0][26] = 8'hd1;
frames[3][0][27] = 8'hd1;
frames[3][0][28] = 8'hd1;
frames[3][0][29] = 8'hd1;
frames[3][0][30] = 8'hd1;
frames[3][0][31] = 8'hd1;
frames[3][0][32] = 8'hd1;
frames[3][0][33] = 8'hd5;
frames[3][0][34] = 8'hd5;
frames[3][0][35] = 8'hd1;
frames[3][0][36] = 8'hd1;
frames[3][0][37] = 8'hd1;
frames[3][0][38] = 8'hb1;
frames[3][0][39] = 8'had;
frames[3][1][0] = 8'hd1;
frames[3][1][1] = 8'hd1;
frames[3][1][2] = 8'hd1;
frames[3][1][3] = 8'hb1;
frames[3][1][4] = 8'hd1;
frames[3][1][5] = 8'hd1;
frames[3][1][6] = 8'hd1;
frames[3][1][7] = 8'hd5;
frames[3][1][8] = 8'hd1;
frames[3][1][9] = 8'hd1;
frames[3][1][10] = 8'hd1;
frames[3][1][11] = 8'hd5;
frames[3][1][12] = 8'hd5;
frames[3][1][13] = 8'hd5;
frames[3][1][14] = 8'hd5;
frames[3][1][15] = 8'hd5;
frames[3][1][16] = 8'hd5;
frames[3][1][17] = 8'hd1;
frames[3][1][18] = 8'hd1;
frames[3][1][19] = 8'hd1;
frames[3][1][20] = 8'hd1;
frames[3][1][21] = 8'hd1;
frames[3][1][22] = 8'hd5;
frames[3][1][23] = 8'hd5;
frames[3][1][24] = 8'hd5;
frames[3][1][25] = 8'hd5;
frames[3][1][26] = 8'hd1;
frames[3][1][27] = 8'hd1;
frames[3][1][28] = 8'hd1;
frames[3][1][29] = 8'hd1;
frames[3][1][30] = 8'hd1;
frames[3][1][31] = 8'hd1;
frames[3][1][32] = 8'hd1;
frames[3][1][33] = 8'hd5;
frames[3][1][34] = 8'hd5;
frames[3][1][35] = 8'hd1;
frames[3][1][36] = 8'hd1;
frames[3][1][37] = 8'hd1;
frames[3][1][38] = 8'hb1;
frames[3][1][39] = 8'had;
frames[3][2][0] = 8'h8d;
frames[3][2][1] = 8'had;
frames[3][2][2] = 8'hd1;
frames[3][2][3] = 8'hd1;
frames[3][2][4] = 8'hd1;
frames[3][2][5] = 8'hd5;
frames[3][2][6] = 8'hf6;
frames[3][2][7] = 8'hd1;
frames[3][2][8] = 8'hd1;
frames[3][2][9] = 8'hd1;
frames[3][2][10] = 8'hd1;
frames[3][2][11] = 8'hd5;
frames[3][2][12] = 8'hd5;
frames[3][2][13] = 8'hd5;
frames[3][2][14] = 8'hd5;
frames[3][2][15] = 8'hd5;
frames[3][2][16] = 8'hd1;
frames[3][2][17] = 8'hd1;
frames[3][2][18] = 8'hd1;
frames[3][2][19] = 8'hd1;
frames[3][2][20] = 8'hd1;
frames[3][2][21] = 8'hd1;
frames[3][2][22] = 8'hd5;
frames[3][2][23] = 8'hd5;
frames[3][2][24] = 8'hd5;
frames[3][2][25] = 8'hd5;
frames[3][2][26] = 8'hd5;
frames[3][2][27] = 8'hd1;
frames[3][2][28] = 8'hd1;
frames[3][2][29] = 8'hd1;
frames[3][2][30] = 8'hd1;
frames[3][2][31] = 8'hd1;
frames[3][2][32] = 8'hd1;
frames[3][2][33] = 8'hd5;
frames[3][2][34] = 8'hd1;
frames[3][2][35] = 8'hd1;
frames[3][2][36] = 8'hd1;
frames[3][2][37] = 8'hd1;
frames[3][2][38] = 8'hb1;
frames[3][2][39] = 8'had;
frames[3][3][0] = 8'h8d;
frames[3][3][1] = 8'h8d;
frames[3][3][2] = 8'had;
frames[3][3][3] = 8'had;
frames[3][3][4] = 8'hb1;
frames[3][3][5] = 8'hd1;
frames[3][3][6] = 8'had;
frames[3][3][7] = 8'had;
frames[3][3][8] = 8'hcd;
frames[3][3][9] = 8'hd1;
frames[3][3][10] = 8'hd1;
frames[3][3][11] = 8'hd5;
frames[3][3][12] = 8'hd5;
frames[3][3][13] = 8'hd5;
frames[3][3][14] = 8'hd5;
frames[3][3][15] = 8'hd5;
frames[3][3][16] = 8'hd1;
frames[3][3][17] = 8'hd1;
frames[3][3][18] = 8'hd1;
frames[3][3][19] = 8'hd1;
frames[3][3][20] = 8'hd1;
frames[3][3][21] = 8'hd1;
frames[3][3][22] = 8'hd5;
frames[3][3][23] = 8'hd5;
frames[3][3][24] = 8'hd5;
frames[3][3][25] = 8'hd5;
frames[3][3][26] = 8'hd5;
frames[3][3][27] = 8'hd1;
frames[3][3][28] = 8'hd1;
frames[3][3][29] = 8'hd1;
frames[3][3][30] = 8'hd1;
frames[3][3][31] = 8'hd1;
frames[3][3][32] = 8'hd1;
frames[3][3][33] = 8'hd5;
frames[3][3][34] = 8'hd1;
frames[3][3][35] = 8'hd1;
frames[3][3][36] = 8'hd1;
frames[3][3][37] = 8'hd1;
frames[3][3][38] = 8'hb1;
frames[3][3][39] = 8'had;
frames[3][4][0] = 8'had;
frames[3][4][1] = 8'had;
frames[3][4][2] = 8'had;
frames[3][4][3] = 8'had;
frames[3][4][4] = 8'had;
frames[3][4][5] = 8'had;
frames[3][4][6] = 8'had;
frames[3][4][7] = 8'h89;
frames[3][4][8] = 8'h84;
frames[3][4][9] = 8'had;
frames[3][4][10] = 8'hd1;
frames[3][4][11] = 8'hd1;
frames[3][4][12] = 8'hd5;
frames[3][4][13] = 8'hd5;
frames[3][4][14] = 8'hd5;
frames[3][4][15] = 8'hd5;
frames[3][4][16] = 8'hd5;
frames[3][4][17] = 8'hd1;
frames[3][4][18] = 8'hd1;
frames[3][4][19] = 8'hd1;
frames[3][4][20] = 8'hd1;
frames[3][4][21] = 8'hd1;
frames[3][4][22] = 8'hd5;
frames[3][4][23] = 8'hd1;
frames[3][4][24] = 8'hd1;
frames[3][4][25] = 8'hd1;
frames[3][4][26] = 8'hd5;
frames[3][4][27] = 8'hd5;
frames[3][4][28] = 8'hd1;
frames[3][4][29] = 8'hd1;
frames[3][4][30] = 8'hd1;
frames[3][4][31] = 8'hd1;
frames[3][4][32] = 8'hd1;
frames[3][4][33] = 8'hd5;
frames[3][4][34] = 8'hd5;
frames[3][4][35] = 8'hd1;
frames[3][4][36] = 8'hd1;
frames[3][4][37] = 8'hd1;
frames[3][4][38] = 8'hd1;
frames[3][4][39] = 8'had;
frames[3][5][0] = 8'had;
frames[3][5][1] = 8'had;
frames[3][5][2] = 8'hb1;
frames[3][5][3] = 8'had;
frames[3][5][4] = 8'had;
frames[3][5][5] = 8'had;
frames[3][5][6] = 8'had;
frames[3][5][7] = 8'had;
frames[3][5][8] = 8'h88;
frames[3][5][9] = 8'h88;
frames[3][5][10] = 8'hb1;
frames[3][5][11] = 8'hd1;
frames[3][5][12] = 8'hd5;
frames[3][5][13] = 8'hd5;
frames[3][5][14] = 8'hd1;
frames[3][5][15] = 8'hd5;
frames[3][5][16] = 8'hd1;
frames[3][5][17] = 8'hb1;
frames[3][5][18] = 8'hd1;
frames[3][5][19] = 8'hd1;
frames[3][5][20] = 8'hb1;
frames[3][5][21] = 8'hb1;
frames[3][5][22] = 8'hd1;
frames[3][5][23] = 8'hd1;
frames[3][5][24] = 8'hd1;
frames[3][5][25] = 8'hd1;
frames[3][5][26] = 8'hd1;
frames[3][5][27] = 8'hd5;
frames[3][5][28] = 8'hd5;
frames[3][5][29] = 8'hd1;
frames[3][5][30] = 8'hd5;
frames[3][5][31] = 8'hd5;
frames[3][5][32] = 8'hd5;
frames[3][5][33] = 8'hd5;
frames[3][5][34] = 8'hd5;
frames[3][5][35] = 8'hd5;
frames[3][5][36] = 8'hd1;
frames[3][5][37] = 8'hd1;
frames[3][5][38] = 8'hd1;
frames[3][5][39] = 8'had;
frames[3][6][0] = 8'hac;
frames[3][6][1] = 8'hac;
frames[3][6][2] = 8'hac;
frames[3][6][3] = 8'hb1;
frames[3][6][4] = 8'hb1;
frames[3][6][5] = 8'hb1;
frames[3][6][6] = 8'had;
frames[3][6][7] = 8'had;
frames[3][6][8] = 8'had;
frames[3][6][9] = 8'had;
frames[3][6][10] = 8'hb1;
frames[3][6][11] = 8'hf6;
frames[3][6][12] = 8'hd6;
frames[3][6][13] = 8'hf6;
frames[3][6][14] = 8'hf6;
frames[3][6][15] = 8'hd5;
frames[3][6][16] = 8'hb5;
frames[3][6][17] = 8'hd5;
frames[3][6][18] = 8'hb1;
frames[3][6][19] = 8'h91;
frames[3][6][20] = 8'h8d;
frames[3][6][21] = 8'hb6;
frames[3][6][22] = 8'hb6;
frames[3][6][23] = 8'h96;
frames[3][6][24] = 8'hb6;
frames[3][6][25] = 8'h96;
frames[3][6][26] = 8'h91;
frames[3][6][27] = 8'h6d;
frames[3][6][28] = 8'h68;
frames[3][6][29] = 8'hd1;
frames[3][6][30] = 8'hd5;
frames[3][6][31] = 8'hf6;
frames[3][6][32] = 8'hd6;
frames[3][6][33] = 8'hd6;
frames[3][6][34] = 8'hd6;
frames[3][6][35] = 8'hd5;
frames[3][6][36] = 8'hd1;
frames[3][6][37] = 8'hd1;
frames[3][6][38] = 8'hd1;
frames[3][6][39] = 8'had;
frames[3][7][0] = 8'hac;
frames[3][7][1] = 8'hac;
frames[3][7][2] = 8'hac;
frames[3][7][3] = 8'hac;
frames[3][7][4] = 8'hac;
frames[3][7][5] = 8'hac;
frames[3][7][6] = 8'had;
frames[3][7][7] = 8'hac;
frames[3][7][8] = 8'h88;
frames[3][7][9] = 8'h8c;
frames[3][7][10] = 8'hd5;
frames[3][7][11] = 8'hfa;
frames[3][7][12] = 8'hfe;
frames[3][7][13] = 8'hfe;
frames[3][7][14] = 8'hfe;
frames[3][7][15] = 8'hd6;
frames[3][7][16] = 8'hb1;
frames[3][7][17] = 8'hb1;
frames[3][7][18] = 8'h6d;
frames[3][7][19] = 8'h69;
frames[3][7][20] = 8'h96;
frames[3][7][21] = 8'h96;
frames[3][7][22] = 8'hb6;
frames[3][7][23] = 8'hda;
frames[3][7][24] = 8'hda;
frames[3][7][25] = 8'hb6;
frames[3][7][26] = 8'h96;
frames[3][7][27] = 8'h49;
frames[3][7][28] = 8'h20;
frames[3][7][29] = 8'hb1;
frames[3][7][30] = 8'hd5;
frames[3][7][31] = 8'hd5;
frames[3][7][32] = 8'hd5;
frames[3][7][33] = 8'hd5;
frames[3][7][34] = 8'hd5;
frames[3][7][35] = 8'hd5;
frames[3][7][36] = 8'hd1;
frames[3][7][37] = 8'hd1;
frames[3][7][38] = 8'hd1;
frames[3][7][39] = 8'had;
frames[3][8][0] = 8'hac;
frames[3][8][1] = 8'hac;
frames[3][8][2] = 8'hac;
frames[3][8][3] = 8'had;
frames[3][8][4] = 8'hac;
frames[3][8][5] = 8'hac;
frames[3][8][6] = 8'hb1;
frames[3][8][7] = 8'hac;
frames[3][8][8] = 8'h8c;
frames[3][8][9] = 8'had;
frames[3][8][10] = 8'hda;
frames[3][8][11] = 8'hfa;
frames[3][8][12] = 8'hfa;
frames[3][8][13] = 8'hfa;
frames[3][8][14] = 8'hfa;
frames[3][8][15] = 8'hfa;
frames[3][8][16] = 8'hb2;
frames[3][8][17] = 8'h8d;
frames[3][8][18] = 8'h6d;
frames[3][8][19] = 8'hb6;
frames[3][8][20] = 8'hb6;
frames[3][8][21] = 8'hba;
frames[3][8][22] = 8'hfa;
frames[3][8][23] = 8'hfa;
frames[3][8][24] = 8'hfa;
frames[3][8][25] = 8'hfa;
frames[3][8][26] = 8'hba;
frames[3][8][27] = 8'h92;
frames[3][8][28] = 8'h44;
frames[3][8][29] = 8'hb1;
frames[3][8][30] = 8'hd1;
frames[3][8][31] = 8'hd5;
frames[3][8][32] = 8'hd1;
frames[3][8][33] = 8'hd5;
frames[3][8][34] = 8'hd5;
frames[3][8][35] = 8'hd5;
frames[3][8][36] = 8'hd1;
frames[3][8][37] = 8'hd1;
frames[3][8][38] = 8'hd1;
frames[3][8][39] = 8'had;
frames[3][9][0] = 8'hac;
frames[3][9][1] = 8'hac;
frames[3][9][2] = 8'had;
frames[3][9][3] = 8'had;
frames[3][9][4] = 8'hac;
frames[3][9][5] = 8'hac;
frames[3][9][6] = 8'hb1;
frames[3][9][7] = 8'hac;
frames[3][9][8] = 8'h8c;
frames[3][9][9] = 8'h8c;
frames[3][9][10] = 8'hb5;
frames[3][9][11] = 8'hfa;
frames[3][9][12] = 8'hfa;
frames[3][9][13] = 8'hfa;
frames[3][9][14] = 8'hfa;
frames[3][9][15] = 8'hfa;
frames[3][9][16] = 8'hb6;
frames[3][9][17] = 8'h91;
frames[3][9][18] = 8'h92;
frames[3][9][19] = 8'hda;
frames[3][9][20] = 8'hfa;
frames[3][9][21] = 8'hfa;
frames[3][9][22] = 8'hfa;
frames[3][9][23] = 8'hfa;
frames[3][9][24] = 8'hfa;
frames[3][9][25] = 8'hfa;
frames[3][9][26] = 8'hfb;
frames[3][9][27] = 8'hda;
frames[3][9][28] = 8'h91;
frames[3][9][29] = 8'hb1;
frames[3][9][30] = 8'hf5;
frames[3][9][31] = 8'hd1;
frames[3][9][32] = 8'hd1;
frames[3][9][33] = 8'hd5;
frames[3][9][34] = 8'hd5;
frames[3][9][35] = 8'hd5;
frames[3][9][36] = 8'hd1;
frames[3][9][37] = 8'hd1;
frames[3][9][38] = 8'hd1;
frames[3][9][39] = 8'hb1;
frames[3][10][0] = 8'hac;
frames[3][10][1] = 8'hac;
frames[3][10][2] = 8'hac;
frames[3][10][3] = 8'hac;
frames[3][10][4] = 8'hac;
frames[3][10][5] = 8'hac;
frames[3][10][6] = 8'hb1;
frames[3][10][7] = 8'hac;
frames[3][10][8] = 8'h8c;
frames[3][10][9] = 8'h8c;
frames[3][10][10] = 8'hd5;
frames[3][10][11] = 8'hfa;
frames[3][10][12] = 8'hfa;
frames[3][10][13] = 8'hfa;
frames[3][10][14] = 8'hfa;
frames[3][10][15] = 8'hfa;
frames[3][10][16] = 8'hb6;
frames[3][10][17] = 8'h91;
frames[3][10][18] = 8'hd6;
frames[3][10][19] = 8'hfb;
frames[3][10][20] = 8'hfa;
frames[3][10][21] = 8'hfa;
frames[3][10][22] = 8'hfa;
frames[3][10][23] = 8'hfa;
frames[3][10][24] = 8'hfa;
frames[3][10][25] = 8'hfa;
frames[3][10][26] = 8'hfa;
frames[3][10][27] = 8'hfa;
frames[3][10][28] = 8'hd6;
frames[3][10][29] = 8'hb6;
frames[3][10][30] = 8'hd1;
frames[3][10][31] = 8'hd1;
frames[3][10][32] = 8'hd1;
frames[3][10][33] = 8'hd1;
frames[3][10][34] = 8'hd5;
frames[3][10][35] = 8'hd5;
frames[3][10][36] = 8'hd1;
frames[3][10][37] = 8'hd1;
frames[3][10][38] = 8'hd1;
frames[3][10][39] = 8'hb1;
frames[3][11][0] = 8'hac;
frames[3][11][1] = 8'hac;
frames[3][11][2] = 8'hac;
frames[3][11][3] = 8'hac;
frames[3][11][4] = 8'hac;
frames[3][11][5] = 8'hac;
frames[3][11][6] = 8'had;
frames[3][11][7] = 8'h8c;
frames[3][11][8] = 8'h88;
frames[3][11][9] = 8'h88;
frames[3][11][10] = 8'hb1;
frames[3][11][11] = 8'hd6;
frames[3][11][12] = 8'hda;
frames[3][11][13] = 8'hfa;
frames[3][11][14] = 8'hfa;
frames[3][11][15] = 8'hfa;
frames[3][11][16] = 8'hb1;
frames[3][11][17] = 8'hb2;
frames[3][11][18] = 8'hda;
frames[3][11][19] = 8'hfb;
frames[3][11][20] = 8'hfb;
frames[3][11][21] = 8'hfb;
frames[3][11][22] = 8'hfa;
frames[3][11][23] = 8'hfa;
frames[3][11][24] = 8'hfa;
frames[3][11][25] = 8'hfa;
frames[3][11][26] = 8'hfa;
frames[3][11][27] = 8'hfa;
frames[3][11][28] = 8'hda;
frames[3][11][29] = 8'hb6;
frames[3][11][30] = 8'hd1;
frames[3][11][31] = 8'hd1;
frames[3][11][32] = 8'hd1;
frames[3][11][33] = 8'hd1;
frames[3][11][34] = 8'hd5;
frames[3][11][35] = 8'hd5;
frames[3][11][36] = 8'hd1;
frames[3][11][37] = 8'hd1;
frames[3][11][38] = 8'hd1;
frames[3][11][39] = 8'hb1;
frames[3][12][0] = 8'h8c;
frames[3][12][1] = 8'hac;
frames[3][12][2] = 8'had;
frames[3][12][3] = 8'hac;
frames[3][12][4] = 8'hac;
frames[3][12][5] = 8'hac;
frames[3][12][6] = 8'had;
frames[3][12][7] = 8'h8c;
frames[3][12][8] = 8'h88;
frames[3][12][9] = 8'h88;
frames[3][12][10] = 8'h8d;
frames[3][12][11] = 8'hd6;
frames[3][12][12] = 8'hfa;
frames[3][12][13] = 8'hfa;
frames[3][12][14] = 8'hfa;
frames[3][12][15] = 8'hd6;
frames[3][12][16] = 8'hb1;
frames[3][12][17] = 8'hd6;
frames[3][12][18] = 8'hfa;
frames[3][12][19] = 8'hfb;
frames[3][12][20] = 8'hff;
frames[3][12][21] = 8'hfa;
frames[3][12][22] = 8'hfa;
frames[3][12][23] = 8'hfa;
frames[3][12][24] = 8'hfa;
frames[3][12][25] = 8'hfa;
frames[3][12][26] = 8'hfa;
frames[3][12][27] = 8'hfa;
frames[3][12][28] = 8'hfa;
frames[3][12][29] = 8'hd6;
frames[3][12][30] = 8'hd1;
frames[3][12][31] = 8'hd1;
frames[3][12][32] = 8'hd1;
frames[3][12][33] = 8'hd1;
frames[3][12][34] = 8'hd5;
frames[3][12][35] = 8'hd5;
frames[3][12][36] = 8'hd1;
frames[3][12][37] = 8'hd1;
frames[3][12][38] = 8'hd1;
frames[3][12][39] = 8'hb1;
frames[3][13][0] = 8'h8c;
frames[3][13][1] = 8'hac;
frames[3][13][2] = 8'had;
frames[3][13][3] = 8'hac;
frames[3][13][4] = 8'hac;
frames[3][13][5] = 8'hac;
frames[3][13][6] = 8'hac;
frames[3][13][7] = 8'h88;
frames[3][13][8] = 8'h88;
frames[3][13][9] = 8'h88;
frames[3][13][10] = 8'h8d;
frames[3][13][11] = 8'hb1;
frames[3][13][12] = 8'hd6;
frames[3][13][13] = 8'hfa;
frames[3][13][14] = 8'hda;
frames[3][13][15] = 8'hb1;
frames[3][13][16] = 8'h91;
frames[3][13][17] = 8'hb6;
frames[3][13][18] = 8'hfa;
frames[3][13][19] = 8'hfb;
frames[3][13][20] = 8'hff;
frames[3][13][21] = 8'hfa;
frames[3][13][22] = 8'hfa;
frames[3][13][23] = 8'hfa;
frames[3][13][24] = 8'hfa;
frames[3][13][25] = 8'hfa;
frames[3][13][26] = 8'hfa;
frames[3][13][27] = 8'hfa;
frames[3][13][28] = 8'hfb;
frames[3][13][29] = 8'hd6;
frames[3][13][30] = 8'hd1;
frames[3][13][31] = 8'hd1;
frames[3][13][32] = 8'hd1;
frames[3][13][33] = 8'hd1;
frames[3][13][34] = 8'hd5;
frames[3][13][35] = 8'hd5;
frames[3][13][36] = 8'hd1;
frames[3][13][37] = 8'hd1;
frames[3][13][38] = 8'hb1;
frames[3][13][39] = 8'hb1;
frames[3][14][0] = 8'h8c;
frames[3][14][1] = 8'hac;
frames[3][14][2] = 8'hac;
frames[3][14][3] = 8'hac;
frames[3][14][4] = 8'hac;
frames[3][14][5] = 8'hac;
frames[3][14][6] = 8'hac;
frames[3][14][7] = 8'h88;
frames[3][14][8] = 8'h88;
frames[3][14][9] = 8'h68;
frames[3][14][10] = 8'h6d;
frames[3][14][11] = 8'h8d;
frames[3][14][12] = 8'hb1;
frames[3][14][13] = 8'hb1;
frames[3][14][14] = 8'hb1;
frames[3][14][15] = 8'hb1;
frames[3][14][16] = 8'h8d;
frames[3][14][17] = 8'hb1;
frames[3][14][18] = 8'hfa;
frames[3][14][19] = 8'hff;
frames[3][14][20] = 8'hff;
frames[3][14][21] = 8'hfb;
frames[3][14][22] = 8'hfa;
frames[3][14][23] = 8'hfa;
frames[3][14][24] = 8'hfa;
frames[3][14][25] = 8'hfa;
frames[3][14][26] = 8'hfa;
frames[3][14][27] = 8'hfa;
frames[3][14][28] = 8'hfa;
frames[3][14][29] = 8'hd6;
frames[3][14][30] = 8'hd1;
frames[3][14][31] = 8'hd1;
frames[3][14][32] = 8'hd1;
frames[3][14][33] = 8'hd1;
frames[3][14][34] = 8'hd1;
frames[3][14][35] = 8'hd5;
frames[3][14][36] = 8'hd1;
frames[3][14][37] = 8'hd1;
frames[3][14][38] = 8'hb1;
frames[3][14][39] = 8'hb1;
frames[3][15][0] = 8'h8c;
frames[3][15][1] = 8'hac;
frames[3][15][2] = 8'hac;
frames[3][15][3] = 8'hac;
frames[3][15][4] = 8'hac;
frames[3][15][5] = 8'hac;
frames[3][15][6] = 8'hac;
frames[3][15][7] = 8'h88;
frames[3][15][8] = 8'h88;
frames[3][15][9] = 8'h68;
frames[3][15][10] = 8'h89;
frames[3][15][11] = 8'h68;
frames[3][15][12] = 8'h69;
frames[3][15][13] = 8'h89;
frames[3][15][14] = 8'h91;
frames[3][15][15] = 8'hb1;
frames[3][15][16] = 8'h8d;
frames[3][15][17] = 8'h8d;
frames[3][15][18] = 8'hfa;
frames[3][15][19] = 8'hff;
frames[3][15][20] = 8'hfb;
frames[3][15][21] = 8'hfb;
frames[3][15][22] = 8'hfb;
frames[3][15][23] = 8'hfa;
frames[3][15][24] = 8'hfa;
frames[3][15][25] = 8'hfa;
frames[3][15][26] = 8'hfa;
frames[3][15][27] = 8'hfa;
frames[3][15][28] = 8'hda;
frames[3][15][29] = 8'hb6;
frames[3][15][30] = 8'hd1;
frames[3][15][31] = 8'hd1;
frames[3][15][32] = 8'hd1;
frames[3][15][33] = 8'hd1;
frames[3][15][34] = 8'hd1;
frames[3][15][35] = 8'hd1;
frames[3][15][36] = 8'hd1;
frames[3][15][37] = 8'hd1;
frames[3][15][38] = 8'hb1;
frames[3][15][39] = 8'hb1;
frames[3][16][0] = 8'h8c;
frames[3][16][1] = 8'hac;
frames[3][16][2] = 8'hac;
frames[3][16][3] = 8'hac;
frames[3][16][4] = 8'hac;
frames[3][16][5] = 8'hac;
frames[3][16][6] = 8'hac;
frames[3][16][7] = 8'h8c;
frames[3][16][8] = 8'h88;
frames[3][16][9] = 8'h68;
frames[3][16][10] = 8'h89;
frames[3][16][11] = 8'h64;
frames[3][16][12] = 8'h60;
frames[3][16][13] = 8'h64;
frames[3][16][14] = 8'h8d;
frames[3][16][15] = 8'hb1;
frames[3][16][16] = 8'h8d;
frames[3][16][17] = 8'h8d;
frames[3][16][18] = 8'hd6;
frames[3][16][19] = 8'hff;
frames[3][16][20] = 8'hfb;
frames[3][16][21] = 8'hfa;
frames[3][16][22] = 8'hfa;
frames[3][16][23] = 8'hfa;
frames[3][16][24] = 8'hfa;
frames[3][16][25] = 8'hfa;
frames[3][16][26] = 8'hfa;
frames[3][16][27] = 8'hfa;
frames[3][16][28] = 8'hda;
frames[3][16][29] = 8'h91;
frames[3][16][30] = 8'hd1;
frames[3][16][31] = 8'hd1;
frames[3][16][32] = 8'hd1;
frames[3][16][33] = 8'hd1;
frames[3][16][34] = 8'hd1;
frames[3][16][35] = 8'hd1;
frames[3][16][36] = 8'hd1;
frames[3][16][37] = 8'hb1;
frames[3][16][38] = 8'hb1;
frames[3][16][39] = 8'hb1;
frames[3][17][0] = 8'h8c;
frames[3][17][1] = 8'hac;
frames[3][17][2] = 8'hac;
frames[3][17][3] = 8'hac;
frames[3][17][4] = 8'hac;
frames[3][17][5] = 8'hac;
frames[3][17][6] = 8'hac;
frames[3][17][7] = 8'h88;
frames[3][17][8] = 8'h68;
frames[3][17][9] = 8'h68;
frames[3][17][10] = 8'h64;
frames[3][17][11] = 8'h40;
frames[3][17][12] = 8'h60;
frames[3][17][13] = 8'h60;
frames[3][17][14] = 8'h69;
frames[3][17][15] = 8'h8d;
frames[3][17][16] = 8'h91;
frames[3][17][17] = 8'h8d;
frames[3][17][18] = 8'hb1;
frames[3][17][19] = 8'hfb;
frames[3][17][20] = 8'hfa;
frames[3][17][21] = 8'hfa;
frames[3][17][22] = 8'hfa;
frames[3][17][23] = 8'hfa;
frames[3][17][24] = 8'hfa;
frames[3][17][25] = 8'hfb;
frames[3][17][26] = 8'hfa;
frames[3][17][27] = 8'hfa;
frames[3][17][28] = 8'hda;
frames[3][17][29] = 8'h6d;
frames[3][17][30] = 8'hb1;
frames[3][17][31] = 8'hd1;
frames[3][17][32] = 8'hd1;
frames[3][17][33] = 8'hd1;
frames[3][17][34] = 8'hd1;
frames[3][17][35] = 8'hd1;
frames[3][17][36] = 8'hd1;
frames[3][17][37] = 8'hb1;
frames[3][17][38] = 8'hb1;
frames[3][17][39] = 8'hb1;
frames[3][18][0] = 8'h8c;
frames[3][18][1] = 8'h8c;
frames[3][18][2] = 8'hac;
frames[3][18][3] = 8'hac;
frames[3][18][4] = 8'hac;
frames[3][18][5] = 8'hac;
frames[3][18][6] = 8'hac;
frames[3][18][7] = 8'hac;
frames[3][18][8] = 8'h88;
frames[3][18][9] = 8'h68;
frames[3][18][10] = 8'h64;
frames[3][18][11] = 8'h40;
frames[3][18][12] = 8'h60;
frames[3][18][13] = 8'h60;
frames[3][18][14] = 8'h69;
frames[3][18][15] = 8'h8d;
frames[3][18][16] = 8'h8d;
frames[3][18][17] = 8'h8d;
frames[3][18][18] = 8'h6d;
frames[3][18][19] = 8'hd6;
frames[3][18][20] = 8'hfa;
frames[3][18][21] = 8'hfa;
frames[3][18][22] = 8'hfa;
frames[3][18][23] = 8'hfa;
frames[3][18][24] = 8'hfa;
frames[3][18][25] = 8'hfa;
frames[3][18][26] = 8'hfa;
frames[3][18][27] = 8'hfa;
frames[3][18][28] = 8'hb6;
frames[3][18][29] = 8'h48;
frames[3][18][30] = 8'hb1;
frames[3][18][31] = 8'hd1;
frames[3][18][32] = 8'hd1;
frames[3][18][33] = 8'hd1;
frames[3][18][34] = 8'hd1;
frames[3][18][35] = 8'hd1;
frames[3][18][36] = 8'hd1;
frames[3][18][37] = 8'hb1;
frames[3][18][38] = 8'hb1;
frames[3][18][39] = 8'hb1;
frames[3][19][0] = 8'h8c;
frames[3][19][1] = 8'h8c;
frames[3][19][2] = 8'hac;
frames[3][19][3] = 8'hac;
frames[3][19][4] = 8'hac;
frames[3][19][5] = 8'hac;
frames[3][19][6] = 8'had;
frames[3][19][7] = 8'hac;
frames[3][19][8] = 8'h88;
frames[3][19][9] = 8'h68;
frames[3][19][10] = 8'h64;
frames[3][19][11] = 8'h40;
frames[3][19][12] = 8'h60;
frames[3][19][13] = 8'h60;
frames[3][19][14] = 8'h68;
frames[3][19][15] = 8'h8d;
frames[3][19][16] = 8'h8d;
frames[3][19][17] = 8'h69;
frames[3][19][18] = 8'h69;
frames[3][19][19] = 8'h8d;
frames[3][19][20] = 8'hda;
frames[3][19][21] = 8'hdb;
frames[3][19][22] = 8'hda;
frames[3][19][23] = 8'hda;
frames[3][19][24] = 8'hda;
frames[3][19][25] = 8'hfa;
frames[3][19][26] = 8'hda;
frames[3][19][27] = 8'hd6;
frames[3][19][28] = 8'h91;
frames[3][19][29] = 8'h44;
frames[3][19][30] = 8'hb1;
frames[3][19][31] = 8'hd1;
frames[3][19][32] = 8'hd1;
frames[3][19][33] = 8'hd1;
frames[3][19][34] = 8'hd1;
frames[3][19][35] = 8'hd1;
frames[3][19][36] = 8'hd1;
frames[3][19][37] = 8'hb1;
frames[3][19][38] = 8'hb1;
frames[3][19][39] = 8'hb1;
frames[3][20][0] = 8'h8c;
frames[3][20][1] = 8'h8c;
frames[3][20][2] = 8'h8c;
frames[3][20][3] = 8'h8c;
frames[3][20][4] = 8'hac;
frames[3][20][5] = 8'hac;
frames[3][20][6] = 8'hac;
frames[3][20][7] = 8'hac;
frames[3][20][8] = 8'h68;
frames[3][20][9] = 8'h88;
frames[3][20][10] = 8'h89;
frames[3][20][11] = 8'h64;
frames[3][20][12] = 8'h64;
frames[3][20][13] = 8'h88;
frames[3][20][14] = 8'h69;
frames[3][20][15] = 8'h8d;
frames[3][20][16] = 8'had;
frames[3][20][17] = 8'h88;
frames[3][20][18] = 8'ha8;
frames[3][20][19] = 8'h84;
frames[3][20][20] = 8'h92;
frames[3][20][21] = 8'hda;
frames[3][20][22] = 8'hb6;
frames[3][20][23] = 8'hb6;
frames[3][20][24] = 8'hb6;
frames[3][20][25] = 8'hda;
frames[3][20][26] = 8'hb6;
frames[3][20][27] = 8'hb6;
frames[3][20][28] = 8'h8d;
frames[3][20][29] = 8'h48;
frames[3][20][30] = 8'hb1;
frames[3][20][31] = 8'hd1;
frames[3][20][32] = 8'hd1;
frames[3][20][33] = 8'hd1;
frames[3][20][34] = 8'hd1;
frames[3][20][35] = 8'hd1;
frames[3][20][36] = 8'hb1;
frames[3][20][37] = 8'hb1;
frames[3][20][38] = 8'hb1;
frames[3][20][39] = 8'hb1;
frames[3][21][0] = 8'h88;
frames[3][21][1] = 8'h88;
frames[3][21][2] = 8'h8c;
frames[3][21][3] = 8'h88;
frames[3][21][4] = 8'h88;
frames[3][21][5] = 8'h8c;
frames[3][21][6] = 8'h8c;
frames[3][21][7] = 8'h8c;
frames[3][21][8] = 8'h68;
frames[3][21][9] = 8'h88;
frames[3][21][10] = 8'h8d;
frames[3][21][11] = 8'h8d;
frames[3][21][12] = 8'h8d;
frames[3][21][13] = 8'h8d;
frames[3][21][14] = 8'h8d;
frames[3][21][15] = 8'h8d;
frames[3][21][16] = 8'ha8;
frames[3][21][17] = 8'h64;
frames[3][21][18] = 8'ha4;
frames[3][21][19] = 8'ha4;
frames[3][21][20] = 8'h8d;
frames[3][21][21] = 8'hb1;
frames[3][21][22] = 8'hb6;
frames[3][21][23] = 8'hb6;
frames[3][21][24] = 8'hb6;
frames[3][21][25] = 8'hb6;
frames[3][21][26] = 8'hb2;
frames[3][21][27] = 8'h91;
frames[3][21][28] = 8'h91;
frames[3][21][29] = 8'h44;
frames[3][21][30] = 8'had;
frames[3][21][31] = 8'hb1;
frames[3][21][32] = 8'hd1;
frames[3][21][33] = 8'hd1;
frames[3][21][34] = 8'hb1;
frames[3][21][35] = 8'hd1;
frames[3][21][36] = 8'hb1;
frames[3][21][37] = 8'hb1;
frames[3][21][38] = 8'hb1;
frames[3][21][39] = 8'hb1;
frames[3][22][0] = 8'h88;
frames[3][22][1] = 8'h88;
frames[3][22][2] = 8'h88;
frames[3][22][3] = 8'h88;
frames[3][22][4] = 8'h88;
frames[3][22][5] = 8'h88;
frames[3][22][6] = 8'h88;
frames[3][22][7] = 8'h88;
frames[3][22][8] = 8'h68;
frames[3][22][9] = 8'h88;
frames[3][22][10] = 8'h8d;
frames[3][22][11] = 8'h8d;
frames[3][22][12] = 8'h8d;
frames[3][22][13] = 8'h6d;
frames[3][22][14] = 8'h8d;
frames[3][22][15] = 8'h8d;
frames[3][22][16] = 8'h88;
frames[3][22][17] = 8'h84;
frames[3][22][18] = 8'ha4;
frames[3][22][19] = 8'ha4;
frames[3][22][20] = 8'h8d;
frames[3][22][21] = 8'had;
frames[3][22][22] = 8'h91;
frames[3][22][23] = 8'h91;
frames[3][22][24] = 8'h91;
frames[3][22][25] = 8'h91;
frames[3][22][26] = 8'h91;
frames[3][22][27] = 8'h91;
frames[3][22][28] = 8'h8d;
frames[3][22][29] = 8'h24;
frames[3][22][30] = 8'h8d;
frames[3][22][31] = 8'hb1;
frames[3][22][32] = 8'hd1;
frames[3][22][33] = 8'hd1;
frames[3][22][34] = 8'hb1;
frames[3][22][35] = 8'hd1;
frames[3][22][36] = 8'hb1;
frames[3][22][37] = 8'hb1;
frames[3][22][38] = 8'hb1;
frames[3][22][39] = 8'hb1;
frames[3][23][0] = 8'h88;
frames[3][23][1] = 8'h88;
frames[3][23][2] = 8'h88;
frames[3][23][3] = 8'h88;
frames[3][23][4] = 8'h88;
frames[3][23][5] = 8'h8c;
frames[3][23][6] = 8'h8c;
frames[3][23][7] = 8'h8c;
frames[3][23][8] = 8'h88;
frames[3][23][9] = 8'h88;
frames[3][23][10] = 8'h68;
frames[3][23][11] = 8'h8d;
frames[3][23][12] = 8'h8d;
frames[3][23][13] = 8'h6d;
frames[3][23][14] = 8'h8d;
frames[3][23][15] = 8'h8d;
frames[3][23][16] = 8'h89;
frames[3][23][17] = 8'h89;
frames[3][23][18] = 8'h84;
frames[3][23][19] = 8'h84;
frames[3][23][20] = 8'h8d;
frames[3][23][21] = 8'h8d;
frames[3][23][22] = 8'h6d;
frames[3][23][23] = 8'h6d;
frames[3][23][24] = 8'h6d;
frames[3][23][25] = 8'h6d;
frames[3][23][26] = 8'h6d;
frames[3][23][27] = 8'h69;
frames[3][23][28] = 8'h44;
frames[3][23][29] = 8'h20;
frames[3][23][30] = 8'had;
frames[3][23][31] = 8'hb1;
frames[3][23][32] = 8'hd1;
frames[3][23][33] = 8'hb1;
frames[3][23][34] = 8'hb1;
frames[3][23][35] = 8'hd1;
frames[3][23][36] = 8'hb1;
frames[3][23][37] = 8'hb1;
frames[3][23][38] = 8'hb1;
frames[3][23][39] = 8'hb1;
frames[3][24][0] = 8'h68;
frames[3][24][1] = 8'h68;
frames[3][24][2] = 8'h88;
frames[3][24][3] = 8'h88;
frames[3][24][4] = 8'had;
frames[3][24][5] = 8'hd1;
frames[3][24][6] = 8'hd1;
frames[3][24][7] = 8'hd1;
frames[3][24][8] = 8'hd1;
frames[3][24][9] = 8'hd1;
frames[3][24][10] = 8'h44;
frames[3][24][11] = 8'h69;
frames[3][24][12] = 8'h69;
frames[3][24][13] = 8'h44;
frames[3][24][14] = 8'h44;
frames[3][24][15] = 8'h68;
frames[3][24][16] = 8'h8d;
frames[3][24][17] = 8'h44;
frames[3][24][18] = 8'h44;
frames[3][24][19] = 8'h68;
frames[3][24][20] = 8'h68;
frames[3][24][21] = 8'h69;
frames[3][24][22] = 8'h69;
frames[3][24][23] = 8'h68;
frames[3][24][24] = 8'h69;
frames[3][24][25] = 8'h69;
frames[3][24][26] = 8'h6d;
frames[3][24][27] = 8'h6d;
frames[3][24][28] = 8'h8d;
frames[3][24][29] = 8'h8d;
frames[3][24][30] = 8'hd1;
frames[3][24][31] = 8'hb1;
frames[3][24][32] = 8'hb1;
frames[3][24][33] = 8'hb1;
frames[3][24][34] = 8'hb1;
frames[3][24][35] = 8'hd1;
frames[3][24][36] = 8'hb1;
frames[3][24][37] = 8'hb1;
frames[3][24][38] = 8'hb1;
frames[3][24][39] = 8'hb1;
frames[3][25][0] = 8'had;
frames[3][25][1] = 8'had;
frames[3][25][2] = 8'hd1;
frames[3][25][3] = 8'hd1;
frames[3][25][4] = 8'hd1;
frames[3][25][5] = 8'hd1;
frames[3][25][6] = 8'hd1;
frames[3][25][7] = 8'had;
frames[3][25][8] = 8'had;
frames[3][25][9] = 8'had;
frames[3][25][10] = 8'h8d;
frames[3][25][11] = 8'hb1;
frames[3][25][12] = 8'h8d;
frames[3][25][13] = 8'h68;
frames[3][25][14] = 8'h8d;
frames[3][25][15] = 8'h8d;
frames[3][25][16] = 8'hd1;
frames[3][25][17] = 8'hb1;
frames[3][25][18] = 8'hb1;
frames[3][25][19] = 8'hb1;
frames[3][25][20] = 8'hb1;
frames[3][25][21] = 8'hd1;
frames[3][25][22] = 8'hd5;
frames[3][25][23] = 8'hd1;
frames[3][25][24] = 8'hd1;
frames[3][25][25] = 8'hd1;
frames[3][25][26] = 8'hd1;
frames[3][25][27] = 8'hd1;
frames[3][25][28] = 8'hd1;
frames[3][25][29] = 8'hd1;
frames[3][25][30] = 8'hb1;
frames[3][25][31] = 8'hb1;
frames[3][25][32] = 8'hb1;
frames[3][25][33] = 8'hb1;
frames[3][25][34] = 8'hb1;
frames[3][25][35] = 8'hb1;
frames[3][25][36] = 8'hb1;
frames[3][25][37] = 8'hb1;
frames[3][25][38] = 8'hb1;
frames[3][25][39] = 8'hb1;
frames[3][26][0] = 8'hd1;
frames[3][26][1] = 8'hb1;
frames[3][26][2] = 8'had;
frames[3][26][3] = 8'had;
frames[3][26][4] = 8'had;
frames[3][26][5] = 8'hd1;
frames[3][26][6] = 8'hd2;
frames[3][26][7] = 8'had;
frames[3][26][8] = 8'ha8;
frames[3][26][9] = 8'had;
frames[3][26][10] = 8'had;
frames[3][26][11] = 8'had;
frames[3][26][12] = 8'hac;
frames[3][26][13] = 8'hb1;
frames[3][26][14] = 8'hb1;
frames[3][26][15] = 8'hb1;
frames[3][26][16] = 8'hb1;
frames[3][26][17] = 8'hb1;
frames[3][26][18] = 8'hb1;
frames[3][26][19] = 8'hd6;
frames[3][26][20] = 8'hd6;
frames[3][26][21] = 8'hd5;
frames[3][26][22] = 8'hd6;
frames[3][26][23] = 8'hd6;
frames[3][26][24] = 8'hd1;
frames[3][26][25] = 8'hd1;
frames[3][26][26] = 8'hd1;
frames[3][26][27] = 8'hb1;
frames[3][26][28] = 8'hb1;
frames[3][26][29] = 8'hb1;
frames[3][26][30] = 8'hb1;
frames[3][26][31] = 8'hb1;
frames[3][26][32] = 8'hb1;
frames[3][26][33] = 8'hb1;
frames[3][26][34] = 8'hb1;
frames[3][26][35] = 8'hb1;
frames[3][26][36] = 8'hb1;
frames[3][26][37] = 8'hb1;
frames[3][26][38] = 8'hb1;
frames[3][26][39] = 8'hb1;
frames[3][27][0] = 8'h8d;
frames[3][27][1] = 8'h8d;
frames[3][27][2] = 8'h8d;
frames[3][27][3] = 8'h89;
frames[3][27][4] = 8'had;
frames[3][27][5] = 8'had;
frames[3][27][6] = 8'had;
frames[3][27][7] = 8'hd1;
frames[3][27][8] = 8'hcd;
frames[3][27][9] = 8'hcd;
frames[3][27][10] = 8'had;
frames[3][27][11] = 8'had;
frames[3][27][12] = 8'hac;
frames[3][27][13] = 8'hb1;
frames[3][27][14] = 8'hb1;
frames[3][27][15] = 8'hb1;
frames[3][27][16] = 8'hac;
frames[3][27][17] = 8'had;
frames[3][27][18] = 8'hb1;
frames[3][27][19] = 8'hd5;
frames[3][27][20] = 8'hd6;
frames[3][27][21] = 8'hd6;
frames[3][27][22] = 8'hd6;
frames[3][27][23] = 8'hd6;
frames[3][27][24] = 8'hd1;
frames[3][27][25] = 8'hb1;
frames[3][27][26] = 8'hd1;
frames[3][27][27] = 8'hb1;
frames[3][27][28] = 8'hb1;
frames[3][27][29] = 8'hb1;
frames[3][27][30] = 8'hb1;
frames[3][27][31] = 8'hb1;
frames[3][27][32] = 8'hb1;
frames[3][27][33] = 8'hb1;
frames[3][27][34] = 8'hb1;
frames[3][27][35] = 8'hb1;
frames[3][27][36] = 8'hb1;
frames[3][27][37] = 8'hb1;
frames[3][27][38] = 8'hb1;
frames[3][27][39] = 8'hb1;
frames[3][28][0] = 8'h88;
frames[3][28][1] = 8'h88;
frames[3][28][2] = 8'h88;
frames[3][28][3] = 8'h88;
frames[3][28][4] = 8'h88;
frames[3][28][5] = 8'h89;
frames[3][28][6] = 8'h89;
frames[3][28][7] = 8'had;
frames[3][28][8] = 8'had;
frames[3][28][9] = 8'hd1;
frames[3][28][10] = 8'hb1;
frames[3][28][11] = 8'had;
frames[3][28][12] = 8'had;
frames[3][28][13] = 8'hb1;
frames[3][28][14] = 8'hb1;
frames[3][28][15] = 8'hb1;
frames[3][28][16] = 8'hac;
frames[3][28][17] = 8'h8c;
frames[3][28][18] = 8'hac;
frames[3][28][19] = 8'had;
frames[3][28][20] = 8'had;
frames[3][28][21] = 8'hb1;
frames[3][28][22] = 8'hd1;
frames[3][28][23] = 8'hd1;
frames[3][28][24] = 8'hd1;
frames[3][28][25] = 8'hd1;
frames[3][28][26] = 8'hd1;
frames[3][28][27] = 8'hb1;
frames[3][28][28] = 8'hb1;
frames[3][28][29] = 8'hb1;
frames[3][28][30] = 8'hb1;
frames[3][28][31] = 8'hb1;
frames[3][28][32] = 8'hb1;
frames[3][28][33] = 8'hb1;
frames[3][28][34] = 8'hb1;
frames[3][28][35] = 8'hb1;
frames[3][28][36] = 8'hb1;
frames[3][28][37] = 8'hb1;
frames[3][28][38] = 8'hb1;
frames[3][28][39] = 8'hb1;
frames[3][29][0] = 8'h68;
frames[3][29][1] = 8'h68;
frames[3][29][2] = 8'h68;
frames[3][29][3] = 8'h68;
frames[3][29][4] = 8'h88;
frames[3][29][5] = 8'h88;
frames[3][29][6] = 8'h89;
frames[3][29][7] = 8'had;
frames[3][29][8] = 8'had;
frames[3][29][9] = 8'had;
frames[3][29][10] = 8'had;
frames[3][29][11] = 8'had;
frames[3][29][12] = 8'hb1;
frames[3][29][13] = 8'hb1;
frames[3][29][14] = 8'hb1;
frames[3][29][15] = 8'hb1;
frames[3][29][16] = 8'hac;
frames[3][29][17] = 8'h8c;
frames[3][29][18] = 8'h8c;
frames[3][29][19] = 8'h8c;
frames[3][29][20] = 8'h8c;
frames[3][29][21] = 8'h8c;
frames[3][29][22] = 8'had;
frames[3][29][23] = 8'hd1;
frames[3][29][24] = 8'hd1;
frames[3][29][25] = 8'hd1;
frames[3][29][26] = 8'hb1;
frames[3][29][27] = 8'hb1;
frames[3][29][28] = 8'hb1;
frames[3][29][29] = 8'hb1;
frames[3][29][30] = 8'hb1;
frames[3][29][31] = 8'hb1;
frames[3][29][32] = 8'hb1;
frames[3][29][33] = 8'hb1;
frames[3][29][34] = 8'hb1;
frames[3][29][35] = 8'hb1;
frames[3][29][36] = 8'hb1;
frames[3][29][37] = 8'hb1;
frames[3][29][38] = 8'hb1;
frames[3][29][39] = 8'hb1;
frames[4][0][0] = 8'hb1;
frames[4][0][1] = 8'hb1;
frames[4][0][2] = 8'hd1;
frames[4][0][3] = 8'hd1;
frames[4][0][4] = 8'hd1;
frames[4][0][5] = 8'hd1;
frames[4][0][6] = 8'hd1;
frames[4][0][7] = 8'hd5;
frames[4][0][8] = 8'hd5;
frames[4][0][9] = 8'hd1;
frames[4][0][10] = 8'hd1;
frames[4][0][11] = 8'hd5;
frames[4][0][12] = 8'hd5;
frames[4][0][13] = 8'hd5;
frames[4][0][14] = 8'hd5;
frames[4][0][15] = 8'hd5;
frames[4][0][16] = 8'hd5;
frames[4][0][17] = 8'hd1;
frames[4][0][18] = 8'hd5;
frames[4][0][19] = 8'hd1;
frames[4][0][20] = 8'hd1;
frames[4][0][21] = 8'hd1;
frames[4][0][22] = 8'hd5;
frames[4][0][23] = 8'hd5;
frames[4][0][24] = 8'hd5;
frames[4][0][25] = 8'hd5;
frames[4][0][26] = 8'hd1;
frames[4][0][27] = 8'hd1;
frames[4][0][28] = 8'hd1;
frames[4][0][29] = 8'hd1;
frames[4][0][30] = 8'hd1;
frames[4][0][31] = 8'hd1;
frames[4][0][32] = 8'hd1;
frames[4][0][33] = 8'hd5;
frames[4][0][34] = 8'hd5;
frames[4][0][35] = 8'hd1;
frames[4][0][36] = 8'hd1;
frames[4][0][37] = 8'hd1;
frames[4][0][38] = 8'hb1;
frames[4][0][39] = 8'had;
frames[4][1][0] = 8'hb1;
frames[4][1][1] = 8'hb1;
frames[4][1][2] = 8'hd1;
frames[4][1][3] = 8'hd1;
frames[4][1][4] = 8'hd1;
frames[4][1][5] = 8'hd1;
frames[4][1][6] = 8'hd1;
frames[4][1][7] = 8'hd5;
frames[4][1][8] = 8'hd1;
frames[4][1][9] = 8'hd1;
frames[4][1][10] = 8'hd1;
frames[4][1][11] = 8'hd5;
frames[4][1][12] = 8'hd5;
frames[4][1][13] = 8'hd5;
frames[4][1][14] = 8'hd5;
frames[4][1][15] = 8'hd5;
frames[4][1][16] = 8'hd5;
frames[4][1][17] = 8'hd1;
frames[4][1][18] = 8'hd1;
frames[4][1][19] = 8'hd1;
frames[4][1][20] = 8'hd1;
frames[4][1][21] = 8'hd1;
frames[4][1][22] = 8'hd5;
frames[4][1][23] = 8'hd5;
frames[4][1][24] = 8'hd5;
frames[4][1][25] = 8'hd5;
frames[4][1][26] = 8'hd1;
frames[4][1][27] = 8'hd1;
frames[4][1][28] = 8'hd1;
frames[4][1][29] = 8'hd1;
frames[4][1][30] = 8'hd1;
frames[4][1][31] = 8'hd1;
frames[4][1][32] = 8'hd1;
frames[4][1][33] = 8'hd5;
frames[4][1][34] = 8'hd5;
frames[4][1][35] = 8'hd1;
frames[4][1][36] = 8'hd1;
frames[4][1][37] = 8'hd1;
frames[4][1][38] = 8'hb1;
frames[4][1][39] = 8'had;
frames[4][2][0] = 8'hb1;
frames[4][2][1] = 8'hb1;
frames[4][2][2] = 8'hd1;
frames[4][2][3] = 8'hd1;
frames[4][2][4] = 8'hd1;
frames[4][2][5] = 8'hd1;
frames[4][2][6] = 8'hd5;
frames[4][2][7] = 8'hd5;
frames[4][2][8] = 8'hd5;
frames[4][2][9] = 8'hd5;
frames[4][2][10] = 8'hd5;
frames[4][2][11] = 8'hd5;
frames[4][2][12] = 8'hf5;
frames[4][2][13] = 8'hd5;
frames[4][2][14] = 8'hd5;
frames[4][2][15] = 8'hd5;
frames[4][2][16] = 8'hd5;
frames[4][2][17] = 8'hd1;
frames[4][2][18] = 8'hd1;
frames[4][2][19] = 8'hd1;
frames[4][2][20] = 8'hd1;
frames[4][2][21] = 8'hd1;
frames[4][2][22] = 8'hd5;
frames[4][2][23] = 8'hd5;
frames[4][2][24] = 8'hd5;
frames[4][2][25] = 8'hd5;
frames[4][2][26] = 8'hd5;
frames[4][2][27] = 8'hd1;
frames[4][2][28] = 8'hd1;
frames[4][2][29] = 8'hd1;
frames[4][2][30] = 8'hd1;
frames[4][2][31] = 8'hd1;
frames[4][2][32] = 8'hd1;
frames[4][2][33] = 8'hd5;
frames[4][2][34] = 8'hd1;
frames[4][2][35] = 8'hd1;
frames[4][2][36] = 8'hd1;
frames[4][2][37] = 8'hd1;
frames[4][2][38] = 8'hb1;
frames[4][2][39] = 8'had;
frames[4][3][0] = 8'hb1;
frames[4][3][1] = 8'hb1;
frames[4][3][2] = 8'hd1;
frames[4][3][3] = 8'hd1;
frames[4][3][4] = 8'hd1;
frames[4][3][5] = 8'hd1;
frames[4][3][6] = 8'hd6;
frames[4][3][7] = 8'hd6;
frames[4][3][8] = 8'hd5;
frames[4][3][9] = 8'hd6;
frames[4][3][10] = 8'hd6;
frames[4][3][11] = 8'hd6;
frames[4][3][12] = 8'hf5;
frames[4][3][13] = 8'hd5;
frames[4][3][14] = 8'hd5;
frames[4][3][15] = 8'hd5;
frames[4][3][16] = 8'hd1;
frames[4][3][17] = 8'hd1;
frames[4][3][18] = 8'hd1;
frames[4][3][19] = 8'hd1;
frames[4][3][20] = 8'hd1;
frames[4][3][21] = 8'hd1;
frames[4][3][22] = 8'hd5;
frames[4][3][23] = 8'hd5;
frames[4][3][24] = 8'hd5;
frames[4][3][25] = 8'hd5;
frames[4][3][26] = 8'hd5;
frames[4][3][27] = 8'hd1;
frames[4][3][28] = 8'hd1;
frames[4][3][29] = 8'hd1;
frames[4][3][30] = 8'hd1;
frames[4][3][31] = 8'hd1;
frames[4][3][32] = 8'hd1;
frames[4][3][33] = 8'hd5;
frames[4][3][34] = 8'hd1;
frames[4][3][35] = 8'hd1;
frames[4][3][36] = 8'hd1;
frames[4][3][37] = 8'hd1;
frames[4][3][38] = 8'hb1;
frames[4][3][39] = 8'had;
frames[4][4][0] = 8'hb1;
frames[4][4][1] = 8'hb1;
frames[4][4][2] = 8'hd1;
frames[4][4][3] = 8'hd1;
frames[4][4][4] = 8'hd1;
frames[4][4][5] = 8'hd1;
frames[4][4][6] = 8'hd1;
frames[4][4][7] = 8'hd5;
frames[4][4][8] = 8'hd5;
frames[4][4][9] = 8'hd1;
frames[4][4][10] = 8'hd5;
frames[4][4][11] = 8'hd5;
frames[4][4][12] = 8'hd5;
frames[4][4][13] = 8'hd5;
frames[4][4][14] = 8'hd5;
frames[4][4][15] = 8'hd5;
frames[4][4][16] = 8'hd1;
frames[4][4][17] = 8'hd1;
frames[4][4][18] = 8'hd1;
frames[4][4][19] = 8'hd1;
frames[4][4][20] = 8'hd1;
frames[4][4][21] = 8'hd1;
frames[4][4][22] = 8'hd5;
frames[4][4][23] = 8'hd1;
frames[4][4][24] = 8'hd1;
frames[4][4][25] = 8'hd1;
frames[4][4][26] = 8'hd1;
frames[4][4][27] = 8'hd1;
frames[4][4][28] = 8'hd1;
frames[4][4][29] = 8'hd1;
frames[4][4][30] = 8'hd1;
frames[4][4][31] = 8'hd1;
frames[4][4][32] = 8'hd1;
frames[4][4][33] = 8'hd5;
frames[4][4][34] = 8'hd5;
frames[4][4][35] = 8'hd1;
frames[4][4][36] = 8'hd1;
frames[4][4][37] = 8'hd1;
frames[4][4][38] = 8'hd1;
frames[4][4][39] = 8'had;
frames[4][5][0] = 8'hb1;
frames[4][5][1] = 8'hb1;
frames[4][5][2] = 8'hd1;
frames[4][5][3] = 8'hd1;
frames[4][5][4] = 8'hd1;
frames[4][5][5] = 8'hd1;
frames[4][5][6] = 8'hd1;
frames[4][5][7] = 8'hd1;
frames[4][5][8] = 8'hd1;
frames[4][5][9] = 8'hb1;
frames[4][5][10] = 8'hb1;
frames[4][5][11] = 8'hd1;
frames[4][5][12] = 8'hd5;
frames[4][5][13] = 8'hd5;
frames[4][5][14] = 8'hd1;
frames[4][5][15] = 8'hd5;
frames[4][5][16] = 8'hd1;
frames[4][5][17] = 8'hd1;
frames[4][5][18] = 8'hd1;
frames[4][5][19] = 8'hd1;
frames[4][5][20] = 8'hb1;
frames[4][5][21] = 8'hb1;
frames[4][5][22] = 8'hd1;
frames[4][5][23] = 8'hd1;
frames[4][5][24] = 8'hd1;
frames[4][5][25] = 8'hd1;
frames[4][5][26] = 8'hd1;
frames[4][5][27] = 8'hd5;
frames[4][5][28] = 8'hd1;
frames[4][5][29] = 8'hd1;
frames[4][5][30] = 8'hd5;
frames[4][5][31] = 8'hd5;
frames[4][5][32] = 8'hd5;
frames[4][5][33] = 8'hd5;
frames[4][5][34] = 8'hd5;
frames[4][5][35] = 8'hd5;
frames[4][5][36] = 8'hd1;
frames[4][5][37] = 8'hd1;
frames[4][5][38] = 8'hd1;
frames[4][5][39] = 8'had;
frames[4][6][0] = 8'hb1;
frames[4][6][1] = 8'hb1;
frames[4][6][2] = 8'hd1;
frames[4][6][3] = 8'hd1;
frames[4][6][4] = 8'hd1;
frames[4][6][5] = 8'hd1;
frames[4][6][6] = 8'hd1;
frames[4][6][7] = 8'hd1;
frames[4][6][8] = 8'hd1;
frames[4][6][9] = 8'hb1;
frames[4][6][10] = 8'hb1;
frames[4][6][11] = 8'hf6;
frames[4][6][12] = 8'hda;
frames[4][6][13] = 8'hd6;
frames[4][6][14] = 8'hfa;
frames[4][6][15] = 8'hd5;
frames[4][6][16] = 8'hb5;
frames[4][6][17] = 8'hd5;
frames[4][6][18] = 8'hb1;
frames[4][6][19] = 8'h91;
frames[4][6][20] = 8'h8d;
frames[4][6][21] = 8'hb6;
frames[4][6][22] = 8'hb6;
frames[4][6][23] = 8'h96;
frames[4][6][24] = 8'hb6;
frames[4][6][25] = 8'h96;
frames[4][6][26] = 8'h91;
frames[4][6][27] = 8'h6d;
frames[4][6][28] = 8'h68;
frames[4][6][29] = 8'hd1;
frames[4][6][30] = 8'hd5;
frames[4][6][31] = 8'hd6;
frames[4][6][32] = 8'hd6;
frames[4][6][33] = 8'hd6;
frames[4][6][34] = 8'hd6;
frames[4][6][35] = 8'hd6;
frames[4][6][36] = 8'hd1;
frames[4][6][37] = 8'hd1;
frames[4][6][38] = 8'hd1;
frames[4][6][39] = 8'had;
frames[4][7][0] = 8'hb1;
frames[4][7][1] = 8'hb1;
frames[4][7][2] = 8'hd1;
frames[4][7][3] = 8'hd1;
frames[4][7][4] = 8'hd1;
frames[4][7][5] = 8'hd1;
frames[4][7][6] = 8'hd1;
frames[4][7][7] = 8'hd1;
frames[4][7][8] = 8'hd1;
frames[4][7][9] = 8'hb1;
frames[4][7][10] = 8'hd6;
frames[4][7][11] = 8'hfe;
frames[4][7][12] = 8'hfe;
frames[4][7][13] = 8'hfe;
frames[4][7][14] = 8'hfa;
frames[4][7][15] = 8'hd6;
frames[4][7][16] = 8'hb1;
frames[4][7][17] = 8'hb1;
frames[4][7][18] = 8'h6d;
frames[4][7][19] = 8'h69;
frames[4][7][20] = 8'h96;
frames[4][7][21] = 8'h96;
frames[4][7][22] = 8'hb6;
frames[4][7][23] = 8'hda;
frames[4][7][24] = 8'hda;
frames[4][7][25] = 8'hb6;
frames[4][7][26] = 8'h96;
frames[4][7][27] = 8'h49;
frames[4][7][28] = 8'h20;
frames[4][7][29] = 8'hb1;
frames[4][7][30] = 8'hd5;
frames[4][7][31] = 8'hd5;
frames[4][7][32] = 8'hd5;
frames[4][7][33] = 8'hd5;
frames[4][7][34] = 8'hd5;
frames[4][7][35] = 8'hd5;
frames[4][7][36] = 8'hd1;
frames[4][7][37] = 8'hd1;
frames[4][7][38] = 8'hd1;
frames[4][7][39] = 8'had;
frames[4][8][0] = 8'had;
frames[4][8][1] = 8'hb1;
frames[4][8][2] = 8'hb1;
frames[4][8][3] = 8'hb1;
frames[4][8][4] = 8'hb1;
frames[4][8][5] = 8'hb1;
frames[4][8][6] = 8'hd1;
frames[4][8][7] = 8'hd1;
frames[4][8][8] = 8'hd1;
frames[4][8][9] = 8'hd5;
frames[4][8][10] = 8'hfa;
frames[4][8][11] = 8'hfa;
frames[4][8][12] = 8'hfa;
frames[4][8][13] = 8'hfa;
frames[4][8][14] = 8'hfa;
frames[4][8][15] = 8'hfa;
frames[4][8][16] = 8'hb1;
frames[4][8][17] = 8'h8d;
frames[4][8][18] = 8'h6d;
frames[4][8][19] = 8'hb6;
frames[4][8][20] = 8'hb6;
frames[4][8][21] = 8'hda;
frames[4][8][22] = 8'hfa;
frames[4][8][23] = 8'hfa;
frames[4][8][24] = 8'hfa;
frames[4][8][25] = 8'hfa;
frames[4][8][26] = 8'hba;
frames[4][8][27] = 8'h92;
frames[4][8][28] = 8'h44;
frames[4][8][29] = 8'hb1;
frames[4][8][30] = 8'hd1;
frames[4][8][31] = 8'hd5;
frames[4][8][32] = 8'hd1;
frames[4][8][33] = 8'hd5;
frames[4][8][34] = 8'hd5;
frames[4][8][35] = 8'hd5;
frames[4][8][36] = 8'hd1;
frames[4][8][37] = 8'hd1;
frames[4][8][38] = 8'hd1;
frames[4][8][39] = 8'had;
frames[4][9][0] = 8'hac;
frames[4][9][1] = 8'hb1;
frames[4][9][2] = 8'hb1;
frames[4][9][3] = 8'hb1;
frames[4][9][4] = 8'hb1;
frames[4][9][5] = 8'hb1;
frames[4][9][6] = 8'hd1;
frames[4][9][7] = 8'hd1;
frames[4][9][8] = 8'hb1;
frames[4][9][9] = 8'hb1;
frames[4][9][10] = 8'hd6;
frames[4][9][11] = 8'hfa;
frames[4][9][12] = 8'hfa;
frames[4][9][13] = 8'hfa;
frames[4][9][14] = 8'hfa;
frames[4][9][15] = 8'hfa;
frames[4][9][16] = 8'hb6;
frames[4][9][17] = 8'h91;
frames[4][9][18] = 8'h92;
frames[4][9][19] = 8'hda;
frames[4][9][20] = 8'hfa;
frames[4][9][21] = 8'hfa;
frames[4][9][22] = 8'hfa;
frames[4][9][23] = 8'hfa;
frames[4][9][24] = 8'hfa;
frames[4][9][25] = 8'hfa;
frames[4][9][26] = 8'hff;
frames[4][9][27] = 8'hda;
frames[4][9][28] = 8'h91;
frames[4][9][29] = 8'hb2;
frames[4][9][30] = 8'hf5;
frames[4][9][31] = 8'hd1;
frames[4][9][32] = 8'hd1;
frames[4][9][33] = 8'hd5;
frames[4][9][34] = 8'hd5;
frames[4][9][35] = 8'hd5;
frames[4][9][36] = 8'hd1;
frames[4][9][37] = 8'hd1;
frames[4][9][38] = 8'hd1;
frames[4][9][39] = 8'hb1;
frames[4][10][0] = 8'hac;
frames[4][10][1] = 8'had;
frames[4][10][2] = 8'hb1;
frames[4][10][3] = 8'hb1;
frames[4][10][4] = 8'hb1;
frames[4][10][5] = 8'hb1;
frames[4][10][6] = 8'hd1;
frames[4][10][7] = 8'hd1;
frames[4][10][8] = 8'hb1;
frames[4][10][9] = 8'had;
frames[4][10][10] = 8'hd6;
frames[4][10][11] = 8'hfa;
frames[4][10][12] = 8'hfa;
frames[4][10][13] = 8'hfa;
frames[4][10][14] = 8'hfa;
frames[4][10][15] = 8'hfa;
frames[4][10][16] = 8'hb6;
frames[4][10][17] = 8'h91;
frames[4][10][18] = 8'hd6;
frames[4][10][19] = 8'hfb;
frames[4][10][20] = 8'hfa;
frames[4][10][21] = 8'hfa;
frames[4][10][22] = 8'hfa;
frames[4][10][23] = 8'hfa;
frames[4][10][24] = 8'hfa;
frames[4][10][25] = 8'hfa;
frames[4][10][26] = 8'hfb;
frames[4][10][27] = 8'hfb;
frames[4][10][28] = 8'hda;
frames[4][10][29] = 8'hb6;
frames[4][10][30] = 8'hd1;
frames[4][10][31] = 8'hd1;
frames[4][10][32] = 8'hd1;
frames[4][10][33] = 8'hd1;
frames[4][10][34] = 8'hd5;
frames[4][10][35] = 8'hd5;
frames[4][10][36] = 8'hd1;
frames[4][10][37] = 8'hd1;
frames[4][10][38] = 8'hd1;
frames[4][10][39] = 8'hb1;
frames[4][11][0] = 8'hac;
frames[4][11][1] = 8'had;
frames[4][11][2] = 8'hb1;
frames[4][11][3] = 8'had;
frames[4][11][4] = 8'hb1;
frames[4][11][5] = 8'hd1;
frames[4][11][6] = 8'hd1;
frames[4][11][7] = 8'hd1;
frames[4][11][8] = 8'hb1;
frames[4][11][9] = 8'hac;
frames[4][11][10] = 8'hd5;
frames[4][11][11] = 8'hda;
frames[4][11][12] = 8'hda;
frames[4][11][13] = 8'hfa;
frames[4][11][14] = 8'hfa;
frames[4][11][15] = 8'hfa;
frames[4][11][16] = 8'hb1;
frames[4][11][17] = 8'hb2;
frames[4][11][18] = 8'hfa;
frames[4][11][19] = 8'hff;
frames[4][11][20] = 8'hfb;
frames[4][11][21] = 8'hfa;
frames[4][11][22] = 8'hfa;
frames[4][11][23] = 8'hfa;
frames[4][11][24] = 8'hfa;
frames[4][11][25] = 8'hfa;
frames[4][11][26] = 8'hfa;
frames[4][11][27] = 8'hfa;
frames[4][11][28] = 8'hda;
frames[4][11][29] = 8'hb6;
frames[4][11][30] = 8'hd1;
frames[4][11][31] = 8'hd1;
frames[4][11][32] = 8'hd1;
frames[4][11][33] = 8'hd1;
frames[4][11][34] = 8'hd5;
frames[4][11][35] = 8'hd5;
frames[4][11][36] = 8'hd1;
frames[4][11][37] = 8'hd1;
frames[4][11][38] = 8'hd1;
frames[4][11][39] = 8'hb1;
frames[4][12][0] = 8'hac;
frames[4][12][1] = 8'hac;
frames[4][12][2] = 8'hb1;
frames[4][12][3] = 8'hb1;
frames[4][12][4] = 8'hb1;
frames[4][12][5] = 8'hb1;
frames[4][12][6] = 8'hd1;
frames[4][12][7] = 8'hd1;
frames[4][12][8] = 8'hb1;
frames[4][12][9] = 8'hac;
frames[4][12][10] = 8'h91;
frames[4][12][11] = 8'hd6;
frames[4][12][12] = 8'hfa;
frames[4][12][13] = 8'hfa;
frames[4][12][14] = 8'hfa;
frames[4][12][15] = 8'hd6;
frames[4][12][16] = 8'h91;
frames[4][12][17] = 8'hb6;
frames[4][12][18] = 8'hfa;
frames[4][12][19] = 8'hfb;
frames[4][12][20] = 8'hff;
frames[4][12][21] = 8'hfa;
frames[4][12][22] = 8'hfa;
frames[4][12][23] = 8'hfa;
frames[4][12][24] = 8'hfa;
frames[4][12][25] = 8'hfa;
frames[4][12][26] = 8'hfa;
frames[4][12][27] = 8'hfa;
frames[4][12][28] = 8'hfa;
frames[4][12][29] = 8'hb6;
frames[4][12][30] = 8'hd1;
frames[4][12][31] = 8'hd1;
frames[4][12][32] = 8'hd1;
frames[4][12][33] = 8'hd1;
frames[4][12][34] = 8'hd5;
frames[4][12][35] = 8'hd5;
frames[4][12][36] = 8'hd1;
frames[4][12][37] = 8'hd1;
frames[4][12][38] = 8'hd1;
frames[4][12][39] = 8'hb1;
frames[4][13][0] = 8'hac;
frames[4][13][1] = 8'hac;
frames[4][13][2] = 8'hb1;
frames[4][13][3] = 8'hb1;
frames[4][13][4] = 8'hb1;
frames[4][13][5] = 8'hb1;
frames[4][13][6] = 8'hb1;
frames[4][13][7] = 8'hb1;
frames[4][13][8] = 8'had;
frames[4][13][9] = 8'hac;
frames[4][13][10] = 8'h8d;
frames[4][13][11] = 8'hb1;
frames[4][13][12] = 8'hd6;
frames[4][13][13] = 8'hfa;
frames[4][13][14] = 8'hda;
frames[4][13][15] = 8'hb1;
frames[4][13][16] = 8'h91;
frames[4][13][17] = 8'hb6;
frames[4][13][18] = 8'hfa;
frames[4][13][19] = 8'hfb;
frames[4][13][20] = 8'hff;
frames[4][13][21] = 8'hfa;
frames[4][13][22] = 8'hfa;
frames[4][13][23] = 8'hfa;
frames[4][13][24] = 8'hfa;
frames[4][13][25] = 8'hfa;
frames[4][13][26] = 8'hfa;
frames[4][13][27] = 8'hfa;
frames[4][13][28] = 8'hfb;
frames[4][13][29] = 8'hd6;
frames[4][13][30] = 8'hd1;
frames[4][13][31] = 8'hd1;
frames[4][13][32] = 8'hd1;
frames[4][13][33] = 8'hd1;
frames[4][13][34] = 8'hd5;
frames[4][13][35] = 8'hd5;
frames[4][13][36] = 8'hd1;
frames[4][13][37] = 8'hd1;
frames[4][13][38] = 8'hb1;
frames[4][13][39] = 8'hb1;
frames[4][14][0] = 8'hac;
frames[4][14][1] = 8'hac;
frames[4][14][2] = 8'hb1;
frames[4][14][3] = 8'had;
frames[4][14][4] = 8'hac;
frames[4][14][5] = 8'hb0;
frames[4][14][6] = 8'hb1;
frames[4][14][7] = 8'had;
frames[4][14][8] = 8'had;
frames[4][14][9] = 8'hac;
frames[4][14][10] = 8'h8d;
frames[4][14][11] = 8'h8d;
frames[4][14][12] = 8'hb1;
frames[4][14][13] = 8'hb1;
frames[4][14][14] = 8'h91;
frames[4][14][15] = 8'hb1;
frames[4][14][16] = 8'h91;
frames[4][14][17] = 8'h91;
frames[4][14][18] = 8'hfa;
frames[4][14][19] = 8'hff;
frames[4][14][20] = 8'hff;
frames[4][14][21] = 8'hfa;
frames[4][14][22] = 8'hfa;
frames[4][14][23] = 8'hfa;
frames[4][14][24] = 8'hfa;
frames[4][14][25] = 8'hfa;
frames[4][14][26] = 8'hfa;
frames[4][14][27] = 8'hfa;
frames[4][14][28] = 8'hfa;
frames[4][14][29] = 8'hd6;
frames[4][14][30] = 8'hd1;
frames[4][14][31] = 8'hd1;
frames[4][14][32] = 8'hd1;
frames[4][14][33] = 8'hd1;
frames[4][14][34] = 8'hd1;
frames[4][14][35] = 8'hd5;
frames[4][14][36] = 8'hd1;
frames[4][14][37] = 8'hd1;
frames[4][14][38] = 8'hb1;
frames[4][14][39] = 8'hb1;
frames[4][15][0] = 8'hac;
frames[4][15][1] = 8'hac;
frames[4][15][2] = 8'had;
frames[4][15][3] = 8'had;
frames[4][15][4] = 8'hac;
frames[4][15][5] = 8'hb1;
frames[4][15][6] = 8'hb1;
frames[4][15][7] = 8'had;
frames[4][15][8] = 8'had;
frames[4][15][9] = 8'hac;
frames[4][15][10] = 8'h8d;
frames[4][15][11] = 8'h69;
frames[4][15][12] = 8'h69;
frames[4][15][13] = 8'h8d;
frames[4][15][14] = 8'h91;
frames[4][15][15] = 8'hb1;
frames[4][15][16] = 8'h8d;
frames[4][15][17] = 8'h8d;
frames[4][15][18] = 8'hfa;
frames[4][15][19] = 8'hff;
frames[4][15][20] = 8'hfb;
frames[4][15][21] = 8'hfb;
frames[4][15][22] = 8'hfb;
frames[4][15][23] = 8'hfa;
frames[4][15][24] = 8'hfa;
frames[4][15][25] = 8'hfa;
frames[4][15][26] = 8'hfa;
frames[4][15][27] = 8'hfa;
frames[4][15][28] = 8'hda;
frames[4][15][29] = 8'hb6;
frames[4][15][30] = 8'hd1;
frames[4][15][31] = 8'hd1;
frames[4][15][32] = 8'hd1;
frames[4][15][33] = 8'hd1;
frames[4][15][34] = 8'hd1;
frames[4][15][35] = 8'hd5;
frames[4][15][36] = 8'hd1;
frames[4][15][37] = 8'hd1;
frames[4][15][38] = 8'hb1;
frames[4][15][39] = 8'hb1;
frames[4][16][0] = 8'hac;
frames[4][16][1] = 8'hac;
frames[4][16][2] = 8'hac;
frames[4][16][3] = 8'hac;
frames[4][16][4] = 8'hac;
frames[4][16][5] = 8'hb1;
frames[4][16][6] = 8'hb1;
frames[4][16][7] = 8'hac;
frames[4][16][8] = 8'had;
frames[4][16][9] = 8'hac;
frames[4][16][10] = 8'ha9;
frames[4][16][11] = 8'h64;
frames[4][16][12] = 8'h60;
frames[4][16][13] = 8'h64;
frames[4][16][14] = 8'h8d;
frames[4][16][15] = 8'hb1;
frames[4][16][16] = 8'h8d;
frames[4][16][17] = 8'h8d;
frames[4][16][18] = 8'hd6;
frames[4][16][19] = 8'hff;
frames[4][16][20] = 8'hfb;
frames[4][16][21] = 8'hfa;
frames[4][16][22] = 8'hfa;
frames[4][16][23] = 8'hfa;
frames[4][16][24] = 8'hfa;
frames[4][16][25] = 8'hfa;
frames[4][16][26] = 8'hfa;
frames[4][16][27] = 8'hfa;
frames[4][16][28] = 8'hda;
frames[4][16][29] = 8'h91;
frames[4][16][30] = 8'hd1;
frames[4][16][31] = 8'hd1;
frames[4][16][32] = 8'hd1;
frames[4][16][33] = 8'hd1;
frames[4][16][34] = 8'hd1;
frames[4][16][35] = 8'hd5;
frames[4][16][36] = 8'hd1;
frames[4][16][37] = 8'hb1;
frames[4][16][38] = 8'hb1;
frames[4][16][39] = 8'hb1;
frames[4][17][0] = 8'hac;
frames[4][17][1] = 8'hac;
frames[4][17][2] = 8'hac;
frames[4][17][3] = 8'hac;
frames[4][17][4] = 8'hac;
frames[4][17][5] = 8'hb1;
frames[4][17][6] = 8'hb1;
frames[4][17][7] = 8'hac;
frames[4][17][8] = 8'hac;
frames[4][17][9] = 8'h8c;
frames[4][17][10] = 8'h84;
frames[4][17][11] = 8'h60;
frames[4][17][12] = 8'h60;
frames[4][17][13] = 8'h60;
frames[4][17][14] = 8'h69;
frames[4][17][15] = 8'h8d;
frames[4][17][16] = 8'h91;
frames[4][17][17] = 8'h8d;
frames[4][17][18] = 8'hb1;
frames[4][17][19] = 8'hfb;
frames[4][17][20] = 8'hfb;
frames[4][17][21] = 8'hfa;
frames[4][17][22] = 8'hfa;
frames[4][17][23] = 8'hfa;
frames[4][17][24] = 8'hfa;
frames[4][17][25] = 8'hfa;
frames[4][17][26] = 8'hfa;
frames[4][17][27] = 8'hfa;
frames[4][17][28] = 8'hb6;
frames[4][17][29] = 8'h6d;
frames[4][17][30] = 8'hb1;
frames[4][17][31] = 8'hd1;
frames[4][17][32] = 8'hd1;
frames[4][17][33] = 8'hd1;
frames[4][17][34] = 8'hd1;
frames[4][17][35] = 8'hd5;
frames[4][17][36] = 8'hd1;
frames[4][17][37] = 8'hb1;
frames[4][17][38] = 8'hb1;
frames[4][17][39] = 8'hb1;
frames[4][18][0] = 8'hac;
frames[4][18][1] = 8'hac;
frames[4][18][2] = 8'hac;
frames[4][18][3] = 8'hac;
frames[4][18][4] = 8'hb0;
frames[4][18][5] = 8'hd1;
frames[4][18][6] = 8'hd1;
frames[4][18][7] = 8'hb1;
frames[4][18][8] = 8'hac;
frames[4][18][9] = 8'h8c;
frames[4][18][10] = 8'h64;
frames[4][18][11] = 8'h60;
frames[4][18][12] = 8'h60;
frames[4][18][13] = 8'h60;
frames[4][18][14] = 8'h68;
frames[4][18][15] = 8'h8d;
frames[4][18][16] = 8'h8d;
frames[4][18][17] = 8'h8d;
frames[4][18][18] = 8'h6d;
frames[4][18][19] = 8'hd6;
frames[4][18][20] = 8'hfa;
frames[4][18][21] = 8'hfa;
frames[4][18][22] = 8'hfa;
frames[4][18][23] = 8'hfa;
frames[4][18][24] = 8'hfa;
frames[4][18][25] = 8'hfa;
frames[4][18][26] = 8'hfa;
frames[4][18][27] = 8'hfa;
frames[4][18][28] = 8'hb2;
frames[4][18][29] = 8'h48;
frames[4][18][30] = 8'hb1;
frames[4][18][31] = 8'hd1;
frames[4][18][32] = 8'hd1;
frames[4][18][33] = 8'hd1;
frames[4][18][34] = 8'hd1;
frames[4][18][35] = 8'hd1;
frames[4][18][36] = 8'hd1;
frames[4][18][37] = 8'hb1;
frames[4][18][38] = 8'hb1;
frames[4][18][39] = 8'hb1;
frames[4][19][0] = 8'hac;
frames[4][19][1] = 8'hac;
frames[4][19][2] = 8'hac;
frames[4][19][3] = 8'hac;
frames[4][19][4] = 8'hac;
frames[4][19][5] = 8'hd1;
frames[4][19][6] = 8'hd1;
frames[4][19][7] = 8'hd1;
frames[4][19][8] = 8'hac;
frames[4][19][9] = 8'h8c;
frames[4][19][10] = 8'h64;
frames[4][19][11] = 8'h40;
frames[4][19][12] = 8'h60;
frames[4][19][13] = 8'h60;
frames[4][19][14] = 8'h68;
frames[4][19][15] = 8'h8d;
frames[4][19][16] = 8'h8d;
frames[4][19][17] = 8'h69;
frames[4][19][18] = 8'h69;
frames[4][19][19] = 8'h8d;
frames[4][19][20] = 8'hda;
frames[4][19][21] = 8'hdb;
frames[4][19][22] = 8'hda;
frames[4][19][23] = 8'hda;
frames[4][19][24] = 8'hda;
frames[4][19][25] = 8'hda;
frames[4][19][26] = 8'hda;
frames[4][19][27] = 8'hb6;
frames[4][19][28] = 8'h8d;
frames[4][19][29] = 8'h44;
frames[4][19][30] = 8'hb1;
frames[4][19][31] = 8'hb1;
frames[4][19][32] = 8'hd1;
frames[4][19][33] = 8'hd1;
frames[4][19][34] = 8'hd1;
frames[4][19][35] = 8'hd1;
frames[4][19][36] = 8'hd1;
frames[4][19][37] = 8'hb1;
frames[4][19][38] = 8'hb1;
frames[4][19][39] = 8'hb1;
frames[4][20][0] = 8'hac;
frames[4][20][1] = 8'hac;
frames[4][20][2] = 8'hac;
frames[4][20][3] = 8'hac;
frames[4][20][4] = 8'hac;
frames[4][20][5] = 8'hb1;
frames[4][20][6] = 8'hd1;
frames[4][20][7] = 8'hd1;
frames[4][20][8] = 8'hac;
frames[4][20][9] = 8'hac;
frames[4][20][10] = 8'h89;
frames[4][20][11] = 8'h64;
frames[4][20][12] = 8'h64;
frames[4][20][13] = 8'h88;
frames[4][20][14] = 8'h69;
frames[4][20][15] = 8'h8d;
frames[4][20][16] = 8'ha9;
frames[4][20][17] = 8'h88;
frames[4][20][18] = 8'ha8;
frames[4][20][19] = 8'h84;
frames[4][20][20] = 8'h92;
frames[4][20][21] = 8'hda;
frames[4][20][22] = 8'hb6;
frames[4][20][23] = 8'h96;
frames[4][20][24] = 8'hb6;
frames[4][20][25] = 8'hba;
frames[4][20][26] = 8'hb6;
frames[4][20][27] = 8'h96;
frames[4][20][28] = 8'h8d;
frames[4][20][29] = 8'h44;
frames[4][20][30] = 8'hb1;
frames[4][20][31] = 8'hb1;
frames[4][20][32] = 8'hd1;
frames[4][20][33] = 8'hd1;
frames[4][20][34] = 8'hd1;
frames[4][20][35] = 8'hd1;
frames[4][20][36] = 8'hb1;
frames[4][20][37] = 8'hb1;
frames[4][20][38] = 8'hb1;
frames[4][20][39] = 8'hb1;
frames[4][21][0] = 8'hac;
frames[4][21][1] = 8'hac;
frames[4][21][2] = 8'had;
frames[4][21][3] = 8'hd1;
frames[4][21][4] = 8'hd1;
frames[4][21][5] = 8'hd1;
frames[4][21][6] = 8'hd5;
frames[4][21][7] = 8'hd5;
frames[4][21][8] = 8'hb1;
frames[4][21][9] = 8'hb1;
frames[4][21][10] = 8'h8d;
frames[4][21][11] = 8'h8d;
frames[4][21][12] = 8'h8d;
frames[4][21][13] = 8'h8d;
frames[4][21][14] = 8'h8d;
frames[4][21][15] = 8'h8d;
frames[4][21][16] = 8'ha8;
frames[4][21][17] = 8'h64;
frames[4][21][18] = 8'ha8;
frames[4][21][19] = 8'ha4;
frames[4][21][20] = 8'h8d;
frames[4][21][21] = 8'hb1;
frames[4][21][22] = 8'hb6;
frames[4][21][23] = 8'hb6;
frames[4][21][24] = 8'hb6;
frames[4][21][25] = 8'hb6;
frames[4][21][26] = 8'hb2;
frames[4][21][27] = 8'hb1;
frames[4][21][28] = 8'h91;
frames[4][21][29] = 8'h44;
frames[4][21][30] = 8'had;
frames[4][21][31] = 8'hb1;
frames[4][21][32] = 8'hd1;
frames[4][21][33] = 8'hd1;
frames[4][21][34] = 8'hb1;
frames[4][21][35] = 8'hd1;
frames[4][21][36] = 8'hb1;
frames[4][21][37] = 8'hb1;
frames[4][21][38] = 8'hb1;
frames[4][21][39] = 8'hb1;
frames[4][22][0] = 8'hac;
frames[4][22][1] = 8'hac;
frames[4][22][2] = 8'hb1;
frames[4][22][3] = 8'hd5;
frames[4][22][4] = 8'hd5;
frames[4][22][5] = 8'hd5;
frames[4][22][6] = 8'hd5;
frames[4][22][7] = 8'hd5;
frames[4][22][8] = 8'hd5;
frames[4][22][9] = 8'hb1;
frames[4][22][10] = 8'h91;
frames[4][22][11] = 8'h91;
frames[4][22][12] = 8'h8d;
frames[4][22][13] = 8'h6d;
frames[4][22][14] = 8'h8d;
frames[4][22][15] = 8'h8d;
frames[4][22][16] = 8'h88;
frames[4][22][17] = 8'h84;
frames[4][22][18] = 8'ha4;
frames[4][22][19] = 8'ha4;
frames[4][22][20] = 8'h8d;
frames[4][22][21] = 8'had;
frames[4][22][22] = 8'h91;
frames[4][22][23] = 8'h91;
frames[4][22][24] = 8'h91;
frames[4][22][25] = 8'h91;
frames[4][22][26] = 8'h91;
frames[4][22][27] = 8'hb1;
frames[4][22][28] = 8'h8d;
frames[4][22][29] = 8'h24;
frames[4][22][30] = 8'h8d;
frames[4][22][31] = 8'hb1;
frames[4][22][32] = 8'hd1;
frames[4][22][33] = 8'hd1;
frames[4][22][34] = 8'hb1;
frames[4][22][35] = 8'hd1;
frames[4][22][36] = 8'hb1;
frames[4][22][37] = 8'hb1;
frames[4][22][38] = 8'hb1;
frames[4][22][39] = 8'hb1;
frames[4][23][0] = 8'hac;
frames[4][23][1] = 8'hac;
frames[4][23][2] = 8'hac;
frames[4][23][3] = 8'hb1;
frames[4][23][4] = 8'hb1;
frames[4][23][5] = 8'hd1;
frames[4][23][6] = 8'hd1;
frames[4][23][7] = 8'hd1;
frames[4][23][8] = 8'hb1;
frames[4][23][9] = 8'had;
frames[4][23][10] = 8'h68;
frames[4][23][11] = 8'h8d;
frames[4][23][12] = 8'h8d;
frames[4][23][13] = 8'h8d;
frames[4][23][14] = 8'h8d;
frames[4][23][15] = 8'h8d;
frames[4][23][16] = 8'h89;
frames[4][23][17] = 8'h89;
frames[4][23][18] = 8'h84;
frames[4][23][19] = 8'h84;
frames[4][23][20] = 8'h8d;
frames[4][23][21] = 8'h8d;
frames[4][23][22] = 8'h6d;
frames[4][23][23] = 8'h6d;
frames[4][23][24] = 8'h6d;
frames[4][23][25] = 8'h6d;
frames[4][23][26] = 8'h6d;
frames[4][23][27] = 8'h6d;
frames[4][23][28] = 8'h44;
frames[4][23][29] = 8'h00;
frames[4][23][30] = 8'had;
frames[4][23][31] = 8'hb1;
frames[4][23][32] = 8'hd1;
frames[4][23][33] = 8'hb1;
frames[4][23][34] = 8'hb1;
frames[4][23][35] = 8'hd1;
frames[4][23][36] = 8'hb1;
frames[4][23][37] = 8'hb1;
frames[4][23][38] = 8'hb1;
frames[4][23][39] = 8'hb1;
frames[4][24][0] = 8'hac;
frames[4][24][1] = 8'hac;
frames[4][24][2] = 8'hac;
frames[4][24][3] = 8'hac;
frames[4][24][4] = 8'had;
frames[4][24][5] = 8'hb1;
frames[4][24][6] = 8'hd1;
frames[4][24][7] = 8'hd1;
frames[4][24][8] = 8'had;
frames[4][24][9] = 8'hac;
frames[4][24][10] = 8'h20;
frames[4][24][11] = 8'h69;
frames[4][24][12] = 8'h8d;
frames[4][24][13] = 8'h44;
frames[4][24][14] = 8'h44;
frames[4][24][15] = 8'h68;
frames[4][24][16] = 8'h8d;
frames[4][24][17] = 8'h44;
frames[4][24][18] = 8'h44;
frames[4][24][19] = 8'h68;
frames[4][24][20] = 8'h68;
frames[4][24][21] = 8'h69;
frames[4][24][22] = 8'h69;
frames[4][24][23] = 8'h68;
frames[4][24][24] = 8'h69;
frames[4][24][25] = 8'h69;
frames[4][24][26] = 8'h6d;
frames[4][24][27] = 8'h6d;
frames[4][24][28] = 8'h8d;
frames[4][24][29] = 8'h8d;
frames[4][24][30] = 8'hd1;
frames[4][24][31] = 8'hb1;
frames[4][24][32] = 8'hb1;
frames[4][24][33] = 8'hb1;
frames[4][24][34] = 8'hb1;
frames[4][24][35] = 8'hd1;
frames[4][24][36] = 8'hb1;
frames[4][24][37] = 8'hb1;
frames[4][24][38] = 8'hb1;
frames[4][24][39] = 8'hb1;
frames[4][25][0] = 8'hac;
frames[4][25][1] = 8'hac;
frames[4][25][2] = 8'hac;
frames[4][25][3] = 8'hac;
frames[4][25][4] = 8'had;
frames[4][25][5] = 8'hb1;
frames[4][25][6] = 8'hd1;
frames[4][25][7] = 8'hd1;
frames[4][25][8] = 8'hd1;
frames[4][25][9] = 8'hb1;
frames[4][25][10] = 8'h8d;
frames[4][25][11] = 8'hb1;
frames[4][25][12] = 8'h8d;
frames[4][25][13] = 8'h8d;
frames[4][25][14] = 8'h8d;
frames[4][25][15] = 8'h8d;
frames[4][25][16] = 8'hd6;
frames[4][25][17] = 8'hb1;
frames[4][25][18] = 8'hb1;
frames[4][25][19] = 8'hb1;
frames[4][25][20] = 8'hb1;
frames[4][25][21] = 8'hd1;
frames[4][25][22] = 8'hd5;
frames[4][25][23] = 8'hd5;
frames[4][25][24] = 8'hd5;
frames[4][25][25] = 8'hd1;
frames[4][25][26] = 8'hd1;
frames[4][25][27] = 8'hd1;
frames[4][25][28] = 8'hd1;
frames[4][25][29] = 8'hd1;
frames[4][25][30] = 8'hb1;
frames[4][25][31] = 8'hb1;
frames[4][25][32] = 8'hb1;
frames[4][25][33] = 8'hb1;
frames[4][25][34] = 8'hb1;
frames[4][25][35] = 8'hb1;
frames[4][25][36] = 8'hb1;
frames[4][25][37] = 8'hb1;
frames[4][25][38] = 8'hb1;
frames[4][25][39] = 8'hb1;
frames[4][26][0] = 8'h8c;
frames[4][26][1] = 8'hac;
frames[4][26][2] = 8'hac;
frames[4][26][3] = 8'hac;
frames[4][26][4] = 8'hac;
frames[4][26][5] = 8'hb1;
frames[4][26][6] = 8'hd1;
frames[4][26][7] = 8'hd1;
frames[4][26][8] = 8'hd1;
frames[4][26][9] = 8'hd1;
frames[4][26][10] = 8'hb1;
frames[4][26][11] = 8'hac;
frames[4][26][12] = 8'had;
frames[4][26][13] = 8'hb1;
frames[4][26][14] = 8'hb1;
frames[4][26][15] = 8'hb1;
frames[4][26][16] = 8'hb1;
frames[4][26][17] = 8'hd1;
frames[4][26][18] = 8'hb1;
frames[4][26][19] = 8'hd6;
frames[4][26][20] = 8'hd6;
frames[4][26][21] = 8'hd6;
frames[4][26][22] = 8'hd6;
frames[4][26][23] = 8'hd6;
frames[4][26][24] = 8'hd1;
frames[4][26][25] = 8'hd1;
frames[4][26][26] = 8'hd1;
frames[4][26][27] = 8'hb1;
frames[4][26][28] = 8'hb1;
frames[4][26][29] = 8'hb1;
frames[4][26][30] = 8'hb1;
frames[4][26][31] = 8'hb1;
frames[4][26][32] = 8'hb1;
frames[4][26][33] = 8'hb1;
frames[4][26][34] = 8'hb1;
frames[4][26][35] = 8'hb1;
frames[4][26][36] = 8'hb1;
frames[4][26][37] = 8'hb1;
frames[4][26][38] = 8'hb1;
frames[4][26][39] = 8'hb1;
frames[4][27][0] = 8'h88;
frames[4][27][1] = 8'h8c;
frames[4][27][2] = 8'h8c;
frames[4][27][3] = 8'hac;
frames[4][27][4] = 8'hac;
frames[4][27][5] = 8'hb1;
frames[4][27][6] = 8'hd1;
frames[4][27][7] = 8'hd1;
frames[4][27][8] = 8'hd1;
frames[4][27][9] = 8'hd1;
frames[4][27][10] = 8'hb1;
frames[4][27][11] = 8'had;
frames[4][27][12] = 8'had;
frames[4][27][13] = 8'hb1;
frames[4][27][14] = 8'hb1;
frames[4][27][15] = 8'hb1;
frames[4][27][16] = 8'hac;
frames[4][27][17] = 8'hac;
frames[4][27][18] = 8'hb1;
frames[4][27][19] = 8'hd5;
frames[4][27][20] = 8'hd6;
frames[4][27][21] = 8'hd6;
frames[4][27][22] = 8'hda;
frames[4][27][23] = 8'hda;
frames[4][27][24] = 8'hd1;
frames[4][27][25] = 8'hb1;
frames[4][27][26] = 8'hd1;
frames[4][27][27] = 8'hb1;
frames[4][27][28] = 8'hb1;
frames[4][27][29] = 8'hb1;
frames[4][27][30] = 8'hb1;
frames[4][27][31] = 8'hb1;
frames[4][27][32] = 8'hb1;
frames[4][27][33] = 8'hb1;
frames[4][27][34] = 8'hb1;
frames[4][27][35] = 8'hb1;
frames[4][27][36] = 8'hb1;
frames[4][27][37] = 8'hb1;
frames[4][27][38] = 8'hb1;
frames[4][27][39] = 8'hb1;
frames[4][28][0] = 8'h88;
frames[4][28][1] = 8'h8c;
frames[4][28][2] = 8'h8c;
frames[4][28][3] = 8'hac;
frames[4][28][4] = 8'hac;
frames[4][28][5] = 8'had;
frames[4][28][6] = 8'hb1;
frames[4][28][7] = 8'hb1;
frames[4][28][8] = 8'hd1;
frames[4][28][9] = 8'hd1;
frames[4][28][10] = 8'hb1;
frames[4][28][11] = 8'hb1;
frames[4][28][12] = 8'hb1;
frames[4][28][13] = 8'hb1;
frames[4][28][14] = 8'hb1;
frames[4][28][15] = 8'hb1;
frames[4][28][16] = 8'hac;
frames[4][28][17] = 8'h8c;
frames[4][28][18] = 8'had;
frames[4][28][19] = 8'had;
frames[4][28][20] = 8'had;
frames[4][28][21] = 8'hb1;
frames[4][28][22] = 8'hd1;
frames[4][28][23] = 8'hd1;
frames[4][28][24] = 8'hd1;
frames[4][28][25] = 8'hd1;
frames[4][28][26] = 8'hb1;
frames[4][28][27] = 8'hb1;
frames[4][28][28] = 8'hb1;
frames[4][28][29] = 8'hb1;
frames[4][28][30] = 8'hb1;
frames[4][28][31] = 8'hb1;
frames[4][28][32] = 8'hb1;
frames[4][28][33] = 8'hb1;
frames[4][28][34] = 8'hb1;
frames[4][28][35] = 8'hb1;
frames[4][28][36] = 8'hb1;
frames[4][28][37] = 8'hb1;
frames[4][28][38] = 8'hb1;
frames[4][28][39] = 8'hb1;
frames[4][29][0] = 8'h88;
frames[4][29][1] = 8'h8c;
frames[4][29][2] = 8'h88;
frames[4][29][3] = 8'h8c;
frames[4][29][4] = 8'hac;
frames[4][29][5] = 8'hac;
frames[4][29][6] = 8'had;
frames[4][29][7] = 8'hb1;
frames[4][29][8] = 8'hd1;
frames[4][29][9] = 8'hd1;
frames[4][29][10] = 8'hb1;
frames[4][29][11] = 8'hb1;
frames[4][29][12] = 8'had;
frames[4][29][13] = 8'hb1;
frames[4][29][14] = 8'hb1;
frames[4][29][15] = 8'hb1;
frames[4][29][16] = 8'hac;
frames[4][29][17] = 8'h8c;
frames[4][29][18] = 8'h8c;
frames[4][29][19] = 8'h8c;
frames[4][29][20] = 8'h8c;
frames[4][29][21] = 8'h8c;
frames[4][29][22] = 8'had;
frames[4][29][23] = 8'hd1;
frames[4][29][24] = 8'hd1;
frames[4][29][25] = 8'hd1;
frames[4][29][26] = 8'hb1;
frames[4][29][27] = 8'hb1;
frames[4][29][28] = 8'hb1;
frames[4][29][29] = 8'hb1;
frames[4][29][30] = 8'hb1;
frames[4][29][31] = 8'hb1;
frames[4][29][32] = 8'hb1;
frames[4][29][33] = 8'hb1;
frames[4][29][34] = 8'hb1;
frames[4][29][35] = 8'hb1;
frames[4][29][36] = 8'hb1;
frames[4][29][37] = 8'hb1;
frames[4][29][38] = 8'hb1;
frames[4][29][39] = 8'hb1;
frames[5][0][0] = 8'hb1;
frames[5][0][1] = 8'hb1;
frames[5][0][2] = 8'hb1;
frames[5][0][3] = 8'hd1;
frames[5][0][4] = 8'hd1;
frames[5][0][5] = 8'hd1;
frames[5][0][6] = 8'hd1;
frames[5][0][7] = 8'hd5;
frames[5][0][8] = 8'hd1;
frames[5][0][9] = 8'hd1;
frames[5][0][10] = 8'hd1;
frames[5][0][11] = 8'hd5;
frames[5][0][12] = 8'hd5;
frames[5][0][13] = 8'hd5;
frames[5][0][14] = 8'hd5;
frames[5][0][15] = 8'hd5;
frames[5][0][16] = 8'hd5;
frames[5][0][17] = 8'hd1;
frames[5][0][18] = 8'hd5;
frames[5][0][19] = 8'hd1;
frames[5][0][20] = 8'hd1;
frames[5][0][21] = 8'hd1;
frames[5][0][22] = 8'hd5;
frames[5][0][23] = 8'hd5;
frames[5][0][24] = 8'hd5;
frames[5][0][25] = 8'hd5;
frames[5][0][26] = 8'hd1;
frames[5][0][27] = 8'hd1;
frames[5][0][28] = 8'hd1;
frames[5][0][29] = 8'hd1;
frames[5][0][30] = 8'hd1;
frames[5][0][31] = 8'hd1;
frames[5][0][32] = 8'hd1;
frames[5][0][33] = 8'hd5;
frames[5][0][34] = 8'hd5;
frames[5][0][35] = 8'hd1;
frames[5][0][36] = 8'hd1;
frames[5][0][37] = 8'hd1;
frames[5][0][38] = 8'hb1;
frames[5][0][39] = 8'had;
frames[5][1][0] = 8'hb1;
frames[5][1][1] = 8'hb1;
frames[5][1][2] = 8'hb1;
frames[5][1][3] = 8'hd1;
frames[5][1][4] = 8'hd1;
frames[5][1][5] = 8'hd1;
frames[5][1][6] = 8'hd1;
frames[5][1][7] = 8'hd1;
frames[5][1][8] = 8'hd1;
frames[5][1][9] = 8'hd1;
frames[5][1][10] = 8'hd1;
frames[5][1][11] = 8'hd5;
frames[5][1][12] = 8'hd5;
frames[5][1][13] = 8'hd5;
frames[5][1][14] = 8'hd5;
frames[5][1][15] = 8'hd5;
frames[5][1][16] = 8'hd5;
frames[5][1][17] = 8'hd1;
frames[5][1][18] = 8'hd1;
frames[5][1][19] = 8'hd1;
frames[5][1][20] = 8'hd1;
frames[5][1][21] = 8'hd1;
frames[5][1][22] = 8'hd5;
frames[5][1][23] = 8'hd5;
frames[5][1][24] = 8'hd5;
frames[5][1][25] = 8'hd5;
frames[5][1][26] = 8'hd1;
frames[5][1][27] = 8'hd1;
frames[5][1][28] = 8'hd1;
frames[5][1][29] = 8'hd1;
frames[5][1][30] = 8'hd1;
frames[5][1][31] = 8'hd1;
frames[5][1][32] = 8'hd1;
frames[5][1][33] = 8'hd5;
frames[5][1][34] = 8'hd5;
frames[5][1][35] = 8'hd1;
frames[5][1][36] = 8'hd1;
frames[5][1][37] = 8'hd1;
frames[5][1][38] = 8'hb1;
frames[5][1][39] = 8'had;
frames[5][2][0] = 8'hb1;
frames[5][2][1] = 8'hb1;
frames[5][2][2] = 8'hd1;
frames[5][2][3] = 8'hd1;
frames[5][2][4] = 8'hd1;
frames[5][2][5] = 8'hd1;
frames[5][2][6] = 8'hd5;
frames[5][2][7] = 8'hd5;
frames[5][2][8] = 8'hd5;
frames[5][2][9] = 8'hd5;
frames[5][2][10] = 8'hd5;
frames[5][2][11] = 8'hd5;
frames[5][2][12] = 8'hf5;
frames[5][2][13] = 8'hd5;
frames[5][2][14] = 8'hd5;
frames[5][2][15] = 8'hd5;
frames[5][2][16] = 8'hd1;
frames[5][2][17] = 8'hd1;
frames[5][2][18] = 8'hd1;
frames[5][2][19] = 8'hd1;
frames[5][2][20] = 8'hd1;
frames[5][2][21] = 8'hd1;
frames[5][2][22] = 8'hd5;
frames[5][2][23] = 8'hd5;
frames[5][2][24] = 8'hd5;
frames[5][2][25] = 8'hd5;
frames[5][2][26] = 8'hd5;
frames[5][2][27] = 8'hd1;
frames[5][2][28] = 8'hd1;
frames[5][2][29] = 8'hd1;
frames[5][2][30] = 8'hd1;
frames[5][2][31] = 8'hd1;
frames[5][2][32] = 8'hd1;
frames[5][2][33] = 8'hd1;
frames[5][2][34] = 8'hd1;
frames[5][2][35] = 8'hd1;
frames[5][2][36] = 8'hd1;
frames[5][2][37] = 8'hd1;
frames[5][2][38] = 8'hb1;
frames[5][2][39] = 8'hac;
frames[5][3][0] = 8'hb1;
frames[5][3][1] = 8'hb1;
frames[5][3][2] = 8'hd1;
frames[5][3][3] = 8'hd1;
frames[5][3][4] = 8'hd1;
frames[5][3][5] = 8'hd1;
frames[5][3][6] = 8'hd6;
frames[5][3][7] = 8'hd6;
frames[5][3][8] = 8'hd6;
frames[5][3][9] = 8'hd6;
frames[5][3][10] = 8'hd6;
frames[5][3][11] = 8'hd6;
frames[5][3][12] = 8'hf6;
frames[5][3][13] = 8'hd5;
frames[5][3][14] = 8'hd5;
frames[5][3][15] = 8'hd5;
frames[5][3][16] = 8'hd1;
frames[5][3][17] = 8'hd1;
frames[5][3][18] = 8'hd1;
frames[5][3][19] = 8'hd1;
frames[5][3][20] = 8'hd1;
frames[5][3][21] = 8'hd1;
frames[5][3][22] = 8'hd5;
frames[5][3][23] = 8'hd5;
frames[5][3][24] = 8'hd5;
frames[5][3][25] = 8'hd5;
frames[5][3][26] = 8'hd5;
frames[5][3][27] = 8'hd1;
frames[5][3][28] = 8'hd1;
frames[5][3][29] = 8'hd1;
frames[5][3][30] = 8'hd1;
frames[5][3][31] = 8'hd1;
frames[5][3][32] = 8'hd1;
frames[5][3][33] = 8'hd5;
frames[5][3][34] = 8'hd1;
frames[5][3][35] = 8'hd1;
frames[5][3][36] = 8'hd1;
frames[5][3][37] = 8'hd1;
frames[5][3][38] = 8'hb1;
frames[5][3][39] = 8'hac;
frames[5][4][0] = 8'hb1;
frames[5][4][1] = 8'hb1;
frames[5][4][2] = 8'hb1;
frames[5][4][3] = 8'hd1;
frames[5][4][4] = 8'hd1;
frames[5][4][5] = 8'hd1;
frames[5][4][6] = 8'hd1;
frames[5][4][7] = 8'hd5;
frames[5][4][8] = 8'hd5;
frames[5][4][9] = 8'hd1;
frames[5][4][10] = 8'hd5;
frames[5][4][11] = 8'hd5;
frames[5][4][12] = 8'hd5;
frames[5][4][13] = 8'hd5;
frames[5][4][14] = 8'hd5;
frames[5][4][15] = 8'hd5;
frames[5][4][16] = 8'hd1;
frames[5][4][17] = 8'hd1;
frames[5][4][18] = 8'hd1;
frames[5][4][19] = 8'hd1;
frames[5][4][20] = 8'hd1;
frames[5][4][21] = 8'hd1;
frames[5][4][22] = 8'hd5;
frames[5][4][23] = 8'hd1;
frames[5][4][24] = 8'hd1;
frames[5][4][25] = 8'hd1;
frames[5][4][26] = 8'hd1;
frames[5][4][27] = 8'hd1;
frames[5][4][28] = 8'hd1;
frames[5][4][29] = 8'hd1;
frames[5][4][30] = 8'hd1;
frames[5][4][31] = 8'hd1;
frames[5][4][32] = 8'hd1;
frames[5][4][33] = 8'hd5;
frames[5][4][34] = 8'hd5;
frames[5][4][35] = 8'hd1;
frames[5][4][36] = 8'hd1;
frames[5][4][37] = 8'hd1;
frames[5][4][38] = 8'hd1;
frames[5][4][39] = 8'had;
frames[5][5][0] = 8'hb1;
frames[5][5][1] = 8'hb1;
frames[5][5][2] = 8'hb1;
frames[5][5][3] = 8'hd1;
frames[5][5][4] = 8'hd1;
frames[5][5][5] = 8'hd1;
frames[5][5][6] = 8'hd1;
frames[5][5][7] = 8'hd1;
frames[5][5][8] = 8'hd1;
frames[5][5][9] = 8'hb1;
frames[5][5][10] = 8'hb1;
frames[5][5][11] = 8'hd1;
frames[5][5][12] = 8'hd5;
frames[5][5][13] = 8'hd5;
frames[5][5][14] = 8'hd1;
frames[5][5][15] = 8'hd5;
frames[5][5][16] = 8'hd1;
frames[5][5][17] = 8'hd1;
frames[5][5][18] = 8'hd1;
frames[5][5][19] = 8'hd1;
frames[5][5][20] = 8'hd1;
frames[5][5][21] = 8'hd1;
frames[5][5][22] = 8'hd1;
frames[5][5][23] = 8'hd1;
frames[5][5][24] = 8'hd1;
frames[5][5][25] = 8'hd1;
frames[5][5][26] = 8'hd1;
frames[5][5][27] = 8'hd1;
frames[5][5][28] = 8'hd1;
frames[5][5][29] = 8'hd1;
frames[5][5][30] = 8'hd5;
frames[5][5][31] = 8'hd5;
frames[5][5][32] = 8'hd5;
frames[5][5][33] = 8'hd5;
frames[5][5][34] = 8'hd5;
frames[5][5][35] = 8'hd5;
frames[5][5][36] = 8'hd1;
frames[5][5][37] = 8'hd1;
frames[5][5][38] = 8'hd1;
frames[5][5][39] = 8'had;
frames[5][6][0] = 8'hb1;
frames[5][6][1] = 8'hb1;
frames[5][6][2] = 8'hd1;
frames[5][6][3] = 8'hd1;
frames[5][6][4] = 8'hd1;
frames[5][6][5] = 8'hd1;
frames[5][6][6] = 8'hd1;
frames[5][6][7] = 8'hd5;
frames[5][6][8] = 8'hd1;
frames[5][6][9] = 8'hb1;
frames[5][6][10] = 8'hd1;
frames[5][6][11] = 8'hfa;
frames[5][6][12] = 8'hda;
frames[5][6][13] = 8'hda;
frames[5][6][14] = 8'hfa;
frames[5][6][15] = 8'hd5;
frames[5][6][16] = 8'hb1;
frames[5][6][17] = 8'hd6;
frames[5][6][18] = 8'hb1;
frames[5][6][19] = 8'hb1;
frames[5][6][20] = 8'h8d;
frames[5][6][21] = 8'hb6;
frames[5][6][22] = 8'hb6;
frames[5][6][23] = 8'h96;
frames[5][6][24] = 8'hb6;
frames[5][6][25] = 8'h96;
frames[5][6][26] = 8'h91;
frames[5][6][27] = 8'h6d;
frames[5][6][28] = 8'h68;
frames[5][6][29] = 8'hd1;
frames[5][6][30] = 8'hd5;
frames[5][6][31] = 8'hd6;
frames[5][6][32] = 8'hd6;
frames[5][6][33] = 8'hd6;
frames[5][6][34] = 8'hd6;
frames[5][6][35] = 8'hd5;
frames[5][6][36] = 8'hd1;
frames[5][6][37] = 8'hd1;
frames[5][6][38] = 8'hd1;
frames[5][6][39] = 8'had;
frames[5][7][0] = 8'hb1;
frames[5][7][1] = 8'hb1;
frames[5][7][2] = 8'hd1;
frames[5][7][3] = 8'hd1;
frames[5][7][4] = 8'hd1;
frames[5][7][5] = 8'hd1;
frames[5][7][6] = 8'hd1;
frames[5][7][7] = 8'hd1;
frames[5][7][8] = 8'hd1;
frames[5][7][9] = 8'hb1;
frames[5][7][10] = 8'hd6;
frames[5][7][11] = 8'hfe;
frames[5][7][12] = 8'hfe;
frames[5][7][13] = 8'hfe;
frames[5][7][14] = 8'hfe;
frames[5][7][15] = 8'hd6;
frames[5][7][16] = 8'hb1;
frames[5][7][17] = 8'hb1;
frames[5][7][18] = 8'h8d;
frames[5][7][19] = 8'h69;
frames[5][7][20] = 8'h96;
frames[5][7][21] = 8'h96;
frames[5][7][22] = 8'hb6;
frames[5][7][23] = 8'hda;
frames[5][7][24] = 8'hda;
frames[5][7][25] = 8'hb6;
frames[5][7][26] = 8'h96;
frames[5][7][27] = 8'h49;
frames[5][7][28] = 8'h20;
frames[5][7][29] = 8'hb1;
frames[5][7][30] = 8'hd5;
frames[5][7][31] = 8'hd5;
frames[5][7][32] = 8'hd5;
frames[5][7][33] = 8'hd5;
frames[5][7][34] = 8'hd5;
frames[5][7][35] = 8'hd5;
frames[5][7][36] = 8'hd1;
frames[5][7][37] = 8'hd1;
frames[5][7][38] = 8'hd1;
frames[5][7][39] = 8'had;
frames[5][8][0] = 8'hac;
frames[5][8][1] = 8'hb1;
frames[5][8][2] = 8'hb1;
frames[5][8][3] = 8'hb1;
frames[5][8][4] = 8'hb1;
frames[5][8][5] = 8'hb1;
frames[5][8][6] = 8'hd1;
frames[5][8][7] = 8'hd1;
frames[5][8][8] = 8'hd1;
frames[5][8][9] = 8'hd5;
frames[5][8][10] = 8'hfa;
frames[5][8][11] = 8'hfa;
frames[5][8][12] = 8'hfa;
frames[5][8][13] = 8'hfa;
frames[5][8][14] = 8'hfa;
frames[5][8][15] = 8'hfa;
frames[5][8][16] = 8'hb1;
frames[5][8][17] = 8'h91;
frames[5][8][18] = 8'h6d;
frames[5][8][19] = 8'hb6;
frames[5][8][20] = 8'hb6;
frames[5][8][21] = 8'hda;
frames[5][8][22] = 8'hfa;
frames[5][8][23] = 8'hfa;
frames[5][8][24] = 8'hfa;
frames[5][8][25] = 8'hfa;
frames[5][8][26] = 8'hba;
frames[5][8][27] = 8'h92;
frames[5][8][28] = 8'h44;
frames[5][8][29] = 8'hb1;
frames[5][8][30] = 8'hd1;
frames[5][8][31] = 8'hd5;
frames[5][8][32] = 8'hd1;
frames[5][8][33] = 8'hd5;
frames[5][8][34] = 8'hd5;
frames[5][8][35] = 8'hd5;
frames[5][8][36] = 8'hd1;
frames[5][8][37] = 8'hd1;
frames[5][8][38] = 8'hd1;
frames[5][8][39] = 8'had;
frames[5][9][0] = 8'hac;
frames[5][9][1] = 8'hb1;
frames[5][9][2] = 8'hb1;
frames[5][9][3] = 8'hb1;
frames[5][9][4] = 8'hb1;
frames[5][9][5] = 8'hb1;
frames[5][9][6] = 8'hd1;
frames[5][9][7] = 8'hd1;
frames[5][9][8] = 8'hb1;
frames[5][9][9] = 8'hb1;
frames[5][9][10] = 8'hd6;
frames[5][9][11] = 8'hfa;
frames[5][9][12] = 8'hfa;
frames[5][9][13] = 8'hfa;
frames[5][9][14] = 8'hfa;
frames[5][9][15] = 8'hfa;
frames[5][9][16] = 8'hb6;
frames[5][9][17] = 8'h91;
frames[5][9][18] = 8'h92;
frames[5][9][19] = 8'hda;
frames[5][9][20] = 8'hfa;
frames[5][9][21] = 8'hfa;
frames[5][9][22] = 8'hfa;
frames[5][9][23] = 8'hfa;
frames[5][9][24] = 8'hfa;
frames[5][9][25] = 8'hfa;
frames[5][9][26] = 8'hff;
frames[5][9][27] = 8'hda;
frames[5][9][28] = 8'h91;
frames[5][9][29] = 8'hb2;
frames[5][9][30] = 8'hf5;
frames[5][9][31] = 8'hd1;
frames[5][9][32] = 8'hd1;
frames[5][9][33] = 8'hd5;
frames[5][9][34] = 8'hd5;
frames[5][9][35] = 8'hd5;
frames[5][9][36] = 8'hd1;
frames[5][9][37] = 8'hd1;
frames[5][9][38] = 8'hd1;
frames[5][9][39] = 8'hb1;
frames[5][10][0] = 8'hac;
frames[5][10][1] = 8'hb1;
frames[5][10][2] = 8'hb1;
frames[5][10][3] = 8'hb1;
frames[5][10][4] = 8'hb1;
frames[5][10][5] = 8'hb1;
frames[5][10][6] = 8'hd1;
frames[5][10][7] = 8'hd1;
frames[5][10][8] = 8'hb1;
frames[5][10][9] = 8'had;
frames[5][10][10] = 8'hd6;
frames[5][10][11] = 8'hfa;
frames[5][10][12] = 8'hfa;
frames[5][10][13] = 8'hfa;
frames[5][10][14] = 8'hfa;
frames[5][10][15] = 8'hfa;
frames[5][10][16] = 8'hb6;
frames[5][10][17] = 8'h91;
frames[5][10][18] = 8'hd6;
frames[5][10][19] = 8'hfb;
frames[5][10][20] = 8'hfa;
frames[5][10][21] = 8'hfa;
frames[5][10][22] = 8'hfa;
frames[5][10][23] = 8'hfa;
frames[5][10][24] = 8'hfa;
frames[5][10][25] = 8'hfa;
frames[5][10][26] = 8'hfb;
frames[5][10][27] = 8'hfb;
frames[5][10][28] = 8'hda;
frames[5][10][29] = 8'hb6;
frames[5][10][30] = 8'hd1;
frames[5][10][31] = 8'hd1;
frames[5][10][32] = 8'hd1;
frames[5][10][33] = 8'hd1;
frames[5][10][34] = 8'hd5;
frames[5][10][35] = 8'hd5;
frames[5][10][36] = 8'hd1;
frames[5][10][37] = 8'hb1;
frames[5][10][38] = 8'hd1;
frames[5][10][39] = 8'hb1;
frames[5][11][0] = 8'hac;
frames[5][11][1] = 8'hac;
frames[5][11][2] = 8'hb1;
frames[5][11][3] = 8'hb1;
frames[5][11][4] = 8'hb1;
frames[5][11][5] = 8'hd1;
frames[5][11][6] = 8'hd1;
frames[5][11][7] = 8'hd1;
frames[5][11][8] = 8'hb1;
frames[5][11][9] = 8'had;
frames[5][11][10] = 8'hd5;
frames[5][11][11] = 8'hda;
frames[5][11][12] = 8'hda;
frames[5][11][13] = 8'hfa;
frames[5][11][14] = 8'hfa;
frames[5][11][15] = 8'hfa;
frames[5][11][16] = 8'hb2;
frames[5][11][17] = 8'hb2;
frames[5][11][18] = 8'hfa;
frames[5][11][19] = 8'hfb;
frames[5][11][20] = 8'hfa;
frames[5][11][21] = 8'hfa;
frames[5][11][22] = 8'hfa;
frames[5][11][23] = 8'hfa;
frames[5][11][24] = 8'hfa;
frames[5][11][25] = 8'hfa;
frames[5][11][26] = 8'hfa;
frames[5][11][27] = 8'hfa;
frames[5][11][28] = 8'hda;
frames[5][11][29] = 8'hb6;
frames[5][11][30] = 8'hd1;
frames[5][11][31] = 8'hd1;
frames[5][11][32] = 8'hd1;
frames[5][11][33] = 8'hd1;
frames[5][11][34] = 8'hd5;
frames[5][11][35] = 8'hd5;
frames[5][11][36] = 8'hd1;
frames[5][11][37] = 8'hb1;
frames[5][11][38] = 8'hd1;
frames[5][11][39] = 8'hb1;
frames[5][12][0] = 8'hac;
frames[5][12][1] = 8'had;
frames[5][12][2] = 8'hb1;
frames[5][12][3] = 8'hb1;
frames[5][12][4] = 8'hb1;
frames[5][12][5] = 8'hb1;
frames[5][12][6] = 8'hd1;
frames[5][12][7] = 8'hb1;
frames[5][12][8] = 8'hb1;
frames[5][12][9] = 8'hac;
frames[5][12][10] = 8'hb1;
frames[5][12][11] = 8'hd6;
frames[5][12][12] = 8'hfa;
frames[5][12][13] = 8'hfa;
frames[5][12][14] = 8'hfa;
frames[5][12][15] = 8'hd6;
frames[5][12][16] = 8'hb1;
frames[5][12][17] = 8'hb6;
frames[5][12][18] = 8'hfa;
frames[5][12][19] = 8'hfb;
frames[5][12][20] = 8'hff;
frames[5][12][21] = 8'hfa;
frames[5][12][22] = 8'hfa;
frames[5][12][23] = 8'hfa;
frames[5][12][24] = 8'hfa;
frames[5][12][25] = 8'hfa;
frames[5][12][26] = 8'hfa;
frames[5][12][27] = 8'hfa;
frames[5][12][28] = 8'hfa;
frames[5][12][29] = 8'hb6;
frames[5][12][30] = 8'hd1;
frames[5][12][31] = 8'hd1;
frames[5][12][32] = 8'hd1;
frames[5][12][33] = 8'hd1;
frames[5][12][34] = 8'hd5;
frames[5][12][35] = 8'hd5;
frames[5][12][36] = 8'hd1;
frames[5][12][37] = 8'hb1;
frames[5][12][38] = 8'hb1;
frames[5][12][39] = 8'hb1;
frames[5][13][0] = 8'hac;
frames[5][13][1] = 8'hac;
frames[5][13][2] = 8'hb1;
frames[5][13][3] = 8'hb1;
frames[5][13][4] = 8'hb1;
frames[5][13][5] = 8'hb1;
frames[5][13][6] = 8'hb1;
frames[5][13][7] = 8'hb1;
frames[5][13][8] = 8'had;
frames[5][13][9] = 8'hac;
frames[5][13][10] = 8'h8d;
frames[5][13][11] = 8'hb1;
frames[5][13][12] = 8'hd6;
frames[5][13][13] = 8'hfa;
frames[5][13][14] = 8'hda;
frames[5][13][15] = 8'hb1;
frames[5][13][16] = 8'h91;
frames[5][13][17] = 8'hb6;
frames[5][13][18] = 8'hfa;
frames[5][13][19] = 8'hff;
frames[5][13][20] = 8'hff;
frames[5][13][21] = 8'hfb;
frames[5][13][22] = 8'hfa;
frames[5][13][23] = 8'hfa;
frames[5][13][24] = 8'hfa;
frames[5][13][25] = 8'hfa;
frames[5][13][26] = 8'hfa;
frames[5][13][27] = 8'hfa;
frames[5][13][28] = 8'hfa;
frames[5][13][29] = 8'hd6;
frames[5][13][30] = 8'hd1;
frames[5][13][31] = 8'hd1;
frames[5][13][32] = 8'hd1;
frames[5][13][33] = 8'hd1;
frames[5][13][34] = 8'hd5;
frames[5][13][35] = 8'hd5;
frames[5][13][36] = 8'hd1;
frames[5][13][37] = 8'hb1;
frames[5][13][38] = 8'hb1;
frames[5][13][39] = 8'hb1;
frames[5][14][0] = 8'hac;
frames[5][14][1] = 8'hac;
frames[5][14][2] = 8'hb1;
frames[5][14][3] = 8'hac;
frames[5][14][4] = 8'hac;
frames[5][14][5] = 8'hb1;
frames[5][14][6] = 8'hb1;
frames[5][14][7] = 8'hac;
frames[5][14][8] = 8'had;
frames[5][14][9] = 8'hac;
frames[5][14][10] = 8'h8d;
frames[5][14][11] = 8'h91;
frames[5][14][12] = 8'hb1;
frames[5][14][13] = 8'hb1;
frames[5][14][14] = 8'h91;
frames[5][14][15] = 8'hb1;
frames[5][14][16] = 8'h91;
frames[5][14][17] = 8'h91;
frames[5][14][18] = 8'hfa;
frames[5][14][19] = 8'hff;
frames[5][14][20] = 8'hff;
frames[5][14][21] = 8'hfa;
frames[5][14][22] = 8'hfa;
frames[5][14][23] = 8'hfa;
frames[5][14][24] = 8'hfa;
frames[5][14][25] = 8'hfa;
frames[5][14][26] = 8'hfa;
frames[5][14][27] = 8'hfa;
frames[5][14][28] = 8'hfa;
frames[5][14][29] = 8'hd6;
frames[5][14][30] = 8'hd1;
frames[5][14][31] = 8'hd1;
frames[5][14][32] = 8'hd1;
frames[5][14][33] = 8'hd1;
frames[5][14][34] = 8'hd5;
frames[5][14][35] = 8'hd5;
frames[5][14][36] = 8'hd1;
frames[5][14][37] = 8'hb1;
frames[5][14][38] = 8'hb1;
frames[5][14][39] = 8'hb1;
frames[5][15][0] = 8'hac;
frames[5][15][1] = 8'hac;
frames[5][15][2] = 8'had;
frames[5][15][3] = 8'had;
frames[5][15][4] = 8'hac;
frames[5][15][5] = 8'hb1;
frames[5][15][6] = 8'hb1;
frames[5][15][7] = 8'hac;
frames[5][15][8] = 8'had;
frames[5][15][9] = 8'hac;
frames[5][15][10] = 8'h8d;
frames[5][15][11] = 8'h68;
frames[5][15][12] = 8'h69;
frames[5][15][13] = 8'h8d;
frames[5][15][14] = 8'h91;
frames[5][15][15] = 8'hb1;
frames[5][15][16] = 8'h8d;
frames[5][15][17] = 8'h8d;
frames[5][15][18] = 8'hfa;
frames[5][15][19] = 8'hff;
frames[5][15][20] = 8'hfb;
frames[5][15][21] = 8'hfb;
frames[5][15][22] = 8'hfa;
frames[5][15][23] = 8'hfa;
frames[5][15][24] = 8'hfa;
frames[5][15][25] = 8'hfa;
frames[5][15][26] = 8'hfa;
frames[5][15][27] = 8'hfa;
frames[5][15][28] = 8'hda;
frames[5][15][29] = 8'hb6;
frames[5][15][30] = 8'hd1;
frames[5][15][31] = 8'hd1;
frames[5][15][32] = 8'hd1;
frames[5][15][33] = 8'hd1;
frames[5][15][34] = 8'hd1;
frames[5][15][35] = 8'hd5;
frames[5][15][36] = 8'hd1;
frames[5][15][37] = 8'hb1;
frames[5][15][38] = 8'hb1;
frames[5][15][39] = 8'hb1;
frames[5][16][0] = 8'hac;
frames[5][16][1] = 8'hac;
frames[5][16][2] = 8'hac;
frames[5][16][3] = 8'hac;
frames[5][16][4] = 8'hac;
frames[5][16][5] = 8'hb1;
frames[5][16][6] = 8'hb1;
frames[5][16][7] = 8'hac;
frames[5][16][8] = 8'hac;
frames[5][16][9] = 8'hac;
frames[5][16][10] = 8'had;
frames[5][16][11] = 8'h64;
frames[5][16][12] = 8'h60;
frames[5][16][13] = 8'h84;
frames[5][16][14] = 8'h8d;
frames[5][16][15] = 8'hb1;
frames[5][16][16] = 8'h8d;
frames[5][16][17] = 8'h8d;
frames[5][16][18] = 8'hd6;
frames[5][16][19] = 8'hff;
frames[5][16][20] = 8'hfa;
frames[5][16][21] = 8'hfa;
frames[5][16][22] = 8'hfa;
frames[5][16][23] = 8'hfa;
frames[5][16][24] = 8'hfa;
frames[5][16][25] = 8'hfa;
frames[5][16][26] = 8'hfa;
frames[5][16][27] = 8'hfa;
frames[5][16][28] = 8'hda;
frames[5][16][29] = 8'h91;
frames[5][16][30] = 8'hb1;
frames[5][16][31] = 8'hd1;
frames[5][16][32] = 8'hd1;
frames[5][16][33] = 8'hd1;
frames[5][16][34] = 8'hd1;
frames[5][16][35] = 8'hd5;
frames[5][16][36] = 8'hd1;
frames[5][16][37] = 8'hb1;
frames[5][16][38] = 8'hb1;
frames[5][16][39] = 8'hb1;
frames[5][17][0] = 8'hac;
frames[5][17][1] = 8'hac;
frames[5][17][2] = 8'hac;
frames[5][17][3] = 8'hac;
frames[5][17][4] = 8'hac;
frames[5][17][5] = 8'hb1;
frames[5][17][6] = 8'hb1;
frames[5][17][7] = 8'hac;
frames[5][17][8] = 8'hac;
frames[5][17][9] = 8'h8c;
frames[5][17][10] = 8'h84;
frames[5][17][11] = 8'h60;
frames[5][17][12] = 8'h60;
frames[5][17][13] = 8'h60;
frames[5][17][14] = 8'h69;
frames[5][17][15] = 8'h8d;
frames[5][17][16] = 8'h91;
frames[5][17][17] = 8'h8d;
frames[5][17][18] = 8'hb1;
frames[5][17][19] = 8'hfb;
frames[5][17][20] = 8'hfa;
frames[5][17][21] = 8'hfa;
frames[5][17][22] = 8'hfa;
frames[5][17][23] = 8'hfa;
frames[5][17][24] = 8'hfa;
frames[5][17][25] = 8'hfa;
frames[5][17][26] = 8'hfa;
frames[5][17][27] = 8'hfa;
frames[5][17][28] = 8'hb6;
frames[5][17][29] = 8'h6d;
frames[5][17][30] = 8'hb1;
frames[5][17][31] = 8'hd1;
frames[5][17][32] = 8'hd1;
frames[5][17][33] = 8'hd1;
frames[5][17][34] = 8'hd1;
frames[5][17][35] = 8'hd1;
frames[5][17][36] = 8'hd1;
frames[5][17][37] = 8'hb1;
frames[5][17][38] = 8'hb1;
frames[5][17][39] = 8'hb1;
frames[5][18][0] = 8'hac;
frames[5][18][1] = 8'hac;
frames[5][18][2] = 8'hac;
frames[5][18][3] = 8'hac;
frames[5][18][4] = 8'hac;
frames[5][18][5] = 8'hd1;
frames[5][18][6] = 8'hd1;
frames[5][18][7] = 8'hb1;
frames[5][18][8] = 8'had;
frames[5][18][9] = 8'h8c;
frames[5][18][10] = 8'h64;
frames[5][18][11] = 8'h60;
frames[5][18][12] = 8'h60;
frames[5][18][13] = 8'h60;
frames[5][18][14] = 8'h68;
frames[5][18][15] = 8'h8d;
frames[5][18][16] = 8'h8d;
frames[5][18][17] = 8'h8d;
frames[5][18][18] = 8'h6d;
frames[5][18][19] = 8'hd6;
frames[5][18][20] = 8'hfa;
frames[5][18][21] = 8'hfa;
frames[5][18][22] = 8'hfa;
frames[5][18][23] = 8'hfa;
frames[5][18][24] = 8'hfa;
frames[5][18][25] = 8'hfa;
frames[5][18][26] = 8'hda;
frames[5][18][27] = 8'hda;
frames[5][18][28] = 8'hb2;
frames[5][18][29] = 8'h48;
frames[5][18][30] = 8'hb1;
frames[5][18][31] = 8'hd1;
frames[5][18][32] = 8'hd1;
frames[5][18][33] = 8'hd1;
frames[5][18][34] = 8'hd1;
frames[5][18][35] = 8'hd1;
frames[5][18][36] = 8'hd1;
frames[5][18][37] = 8'hb1;
frames[5][18][38] = 8'hb1;
frames[5][18][39] = 8'hb1;
frames[5][19][0] = 8'hac;
frames[5][19][1] = 8'hac;
frames[5][19][2] = 8'hac;
frames[5][19][3] = 8'hac;
frames[5][19][4] = 8'hac;
frames[5][19][5] = 8'hd1;
frames[5][19][6] = 8'hd1;
frames[5][19][7] = 8'hd1;
frames[5][19][8] = 8'hac;
frames[5][19][9] = 8'h8c;
frames[5][19][10] = 8'h84;
frames[5][19][11] = 8'h40;
frames[5][19][12] = 8'h60;
frames[5][19][13] = 8'h60;
frames[5][19][14] = 8'h68;
frames[5][19][15] = 8'h8d;
frames[5][19][16] = 8'h8d;
frames[5][19][17] = 8'h69;
frames[5][19][18] = 8'h68;
frames[5][19][19] = 8'h8d;
frames[5][19][20] = 8'hda;
frames[5][19][21] = 8'hdb;
frames[5][19][22] = 8'hfa;
frames[5][19][23] = 8'hda;
frames[5][19][24] = 8'hda;
frames[5][19][25] = 8'hda;
frames[5][19][26] = 8'hda;
frames[5][19][27] = 8'hb6;
frames[5][19][28] = 8'h8d;
frames[5][19][29] = 8'h44;
frames[5][19][30] = 8'hb1;
frames[5][19][31] = 8'hb1;
frames[5][19][32] = 8'hd1;
frames[5][19][33] = 8'hd1;
frames[5][19][34] = 8'hd1;
frames[5][19][35] = 8'hd1;
frames[5][19][36] = 8'hd1;
frames[5][19][37] = 8'hb1;
frames[5][19][38] = 8'hb1;
frames[5][19][39] = 8'hb1;
frames[5][20][0] = 8'hac;
frames[5][20][1] = 8'hac;
frames[5][20][2] = 8'hac;
frames[5][20][3] = 8'hac;
frames[5][20][4] = 8'hac;
frames[5][20][5] = 8'hb1;
frames[5][20][6] = 8'hd1;
frames[5][20][7] = 8'hb1;
frames[5][20][8] = 8'hac;
frames[5][20][9] = 8'hac;
frames[5][20][10] = 8'h89;
frames[5][20][11] = 8'h64;
frames[5][20][12] = 8'h64;
frames[5][20][13] = 8'h88;
frames[5][20][14] = 8'h69;
frames[5][20][15] = 8'h8d;
frames[5][20][16] = 8'ha9;
frames[5][20][17] = 8'h84;
frames[5][20][18] = 8'ha8;
frames[5][20][19] = 8'ha4;
frames[5][20][20] = 8'h92;
frames[5][20][21] = 8'hba;
frames[5][20][22] = 8'hb6;
frames[5][20][23] = 8'h96;
frames[5][20][24] = 8'hb6;
frames[5][20][25] = 8'hba;
frames[5][20][26] = 8'hb6;
frames[5][20][27] = 8'hb6;
frames[5][20][28] = 8'h8d;
frames[5][20][29] = 8'h44;
frames[5][20][30] = 8'hb1;
frames[5][20][31] = 8'hb1;
frames[5][20][32] = 8'hd1;
frames[5][20][33] = 8'hd1;
frames[5][20][34] = 8'hd1;
frames[5][20][35] = 8'hd1;
frames[5][20][36] = 8'hb1;
frames[5][20][37] = 8'hb1;
frames[5][20][38] = 8'hb1;
frames[5][20][39] = 8'hb1;
frames[5][21][0] = 8'hac;
frames[5][21][1] = 8'hac;
frames[5][21][2] = 8'hb1;
frames[5][21][3] = 8'hd1;
frames[5][21][4] = 8'hd1;
frames[5][21][5] = 8'hd1;
frames[5][21][6] = 8'hd5;
frames[5][21][7] = 8'hd5;
frames[5][21][8] = 8'hb1;
frames[5][21][9] = 8'hb1;
frames[5][21][10] = 8'h8d;
frames[5][21][11] = 8'h8d;
frames[5][21][12] = 8'h91;
frames[5][21][13] = 8'h8d;
frames[5][21][14] = 8'h8d;
frames[5][21][15] = 8'h8d;
frames[5][21][16] = 8'ha8;
frames[5][21][17] = 8'h64;
frames[5][21][18] = 8'ha8;
frames[5][21][19] = 8'ha4;
frames[5][21][20] = 8'h8d;
frames[5][21][21] = 8'hb1;
frames[5][21][22] = 8'hb6;
frames[5][21][23] = 8'hb6;
frames[5][21][24] = 8'hb6;
frames[5][21][25] = 8'hb6;
frames[5][21][26] = 8'hb2;
frames[5][21][27] = 8'hb2;
frames[5][21][28] = 8'h91;
frames[5][21][29] = 8'h44;
frames[5][21][30] = 8'had;
frames[5][21][31] = 8'hb1;
frames[5][21][32] = 8'hd1;
frames[5][21][33] = 8'hd1;
frames[5][21][34] = 8'hb1;
frames[5][21][35] = 8'hd1;
frames[5][21][36] = 8'hb1;
frames[5][21][37] = 8'hb1;
frames[5][21][38] = 8'hb1;
frames[5][21][39] = 8'hb1;
frames[5][22][0] = 8'hac;
frames[5][22][1] = 8'hac;
frames[5][22][2] = 8'hb1;
frames[5][22][3] = 8'hd5;
frames[5][22][4] = 8'hd5;
frames[5][22][5] = 8'hd5;
frames[5][22][6] = 8'hd5;
frames[5][22][7] = 8'hd6;
frames[5][22][8] = 8'hb1;
frames[5][22][9] = 8'hb1;
frames[5][22][10] = 8'h91;
frames[5][22][11] = 8'h91;
frames[5][22][12] = 8'h8d;
frames[5][22][13] = 8'h6d;
frames[5][22][14] = 8'h8d;
frames[5][22][15] = 8'h8d;
frames[5][22][16] = 8'h88;
frames[5][22][17] = 8'h84;
frames[5][22][18] = 8'ha4;
frames[5][22][19] = 8'ha8;
frames[5][22][20] = 8'h8d;
frames[5][22][21] = 8'hb1;
frames[5][22][22] = 8'h91;
frames[5][22][23] = 8'h91;
frames[5][22][24] = 8'h91;
frames[5][22][25] = 8'h91;
frames[5][22][26] = 8'h91;
frames[5][22][27] = 8'hb1;
frames[5][22][28] = 8'h8d;
frames[5][22][29] = 8'h24;
frames[5][22][30] = 8'h8d;
frames[5][22][31] = 8'hb1;
frames[5][22][32] = 8'hd1;
frames[5][22][33] = 8'hd1;
frames[5][22][34] = 8'hb1;
frames[5][22][35] = 8'hd1;
frames[5][22][36] = 8'hb1;
frames[5][22][37] = 8'hb1;
frames[5][22][38] = 8'hb1;
frames[5][22][39] = 8'hb1;
frames[5][23][0] = 8'hac;
frames[5][23][1] = 8'hac;
frames[5][23][2] = 8'hac;
frames[5][23][3] = 8'hb1;
frames[5][23][4] = 8'hb1;
frames[5][23][5] = 8'hd1;
frames[5][23][6] = 8'hd1;
frames[5][23][7] = 8'hd1;
frames[5][23][8] = 8'hb1;
frames[5][23][9] = 8'had;
frames[5][23][10] = 8'h68;
frames[5][23][11] = 8'h8d;
frames[5][23][12] = 8'h8d;
frames[5][23][13] = 8'h8d;
frames[5][23][14] = 8'h8d;
frames[5][23][15] = 8'h8d;
frames[5][23][16] = 8'h89;
frames[5][23][17] = 8'h89;
frames[5][23][18] = 8'h84;
frames[5][23][19] = 8'h84;
frames[5][23][20] = 8'h8d;
frames[5][23][21] = 8'h8d;
frames[5][23][22] = 8'h6d;
frames[5][23][23] = 8'h6d;
frames[5][23][24] = 8'h6d;
frames[5][23][25] = 8'h6d;
frames[5][23][26] = 8'h6d;
frames[5][23][27] = 8'h6d;
frames[5][23][28] = 8'h44;
frames[5][23][29] = 8'h00;
frames[5][23][30] = 8'h8d;
frames[5][23][31] = 8'hb1;
frames[5][23][32] = 8'hd1;
frames[5][23][33] = 8'hd1;
frames[5][23][34] = 8'hb1;
frames[5][23][35] = 8'hd1;
frames[5][23][36] = 8'hb1;
frames[5][23][37] = 8'hb1;
frames[5][23][38] = 8'hb1;
frames[5][23][39] = 8'hb1;
frames[5][24][0] = 8'hac;
frames[5][24][1] = 8'hac;
frames[5][24][2] = 8'hac;
frames[5][24][3] = 8'hac;
frames[5][24][4] = 8'hac;
frames[5][24][5] = 8'hd1;
frames[5][24][6] = 8'hd1;
frames[5][24][7] = 8'hd1;
frames[5][24][8] = 8'hb1;
frames[5][24][9] = 8'hac;
frames[5][24][10] = 8'h20;
frames[5][24][11] = 8'h69;
frames[5][24][12] = 8'h8d;
frames[5][24][13] = 8'h44;
frames[5][24][14] = 8'h44;
frames[5][24][15] = 8'h68;
frames[5][24][16] = 8'h8d;
frames[5][24][17] = 8'h44;
frames[5][24][18] = 8'h44;
frames[5][24][19] = 8'h68;
frames[5][24][20] = 8'h68;
frames[5][24][21] = 8'h69;
frames[5][24][22] = 8'h69;
frames[5][24][23] = 8'h69;
frames[5][24][24] = 8'h69;
frames[5][24][25] = 8'h69;
frames[5][24][26] = 8'h6d;
frames[5][24][27] = 8'h6d;
frames[5][24][28] = 8'h6d;
frames[5][24][29] = 8'h8d;
frames[5][24][30] = 8'hd1;
frames[5][24][31] = 8'hb1;
frames[5][24][32] = 8'hb1;
frames[5][24][33] = 8'hb1;
frames[5][24][34] = 8'hb1;
frames[5][24][35] = 8'hb1;
frames[5][24][36] = 8'hb1;
frames[5][24][37] = 8'hb1;
frames[5][24][38] = 8'hb1;
frames[5][24][39] = 8'hb1;
frames[5][25][0] = 8'h8c;
frames[5][25][1] = 8'hac;
frames[5][25][2] = 8'hac;
frames[5][25][3] = 8'hac;
frames[5][25][4] = 8'had;
frames[5][25][5] = 8'hb1;
frames[5][25][6] = 8'hd1;
frames[5][25][7] = 8'hd1;
frames[5][25][8] = 8'hd1;
frames[5][25][9] = 8'hd1;
frames[5][25][10] = 8'h8d;
frames[5][25][11] = 8'hb1;
frames[5][25][12] = 8'h8d;
frames[5][25][13] = 8'h8d;
frames[5][25][14] = 8'h8d;
frames[5][25][15] = 8'h8d;
frames[5][25][16] = 8'hb6;
frames[5][25][17] = 8'h91;
frames[5][25][18] = 8'hb1;
frames[5][25][19] = 8'hb1;
frames[5][25][20] = 8'hb1;
frames[5][25][21] = 8'hb1;
frames[5][25][22] = 8'hd5;
frames[5][25][23] = 8'hd5;
frames[5][25][24] = 8'hd1;
frames[5][25][25] = 8'hd1;
frames[5][25][26] = 8'hd1;
frames[5][25][27] = 8'hd1;
frames[5][25][28] = 8'hd1;
frames[5][25][29] = 8'hd1;
frames[5][25][30] = 8'hb1;
frames[5][25][31] = 8'hb1;
frames[5][25][32] = 8'hb1;
frames[5][25][33] = 8'hb1;
frames[5][25][34] = 8'hb1;
frames[5][25][35] = 8'hb1;
frames[5][25][36] = 8'hb1;
frames[5][25][37] = 8'hb1;
frames[5][25][38] = 8'hb1;
frames[5][25][39] = 8'hb1;
frames[5][26][0] = 8'h8c;
frames[5][26][1] = 8'hac;
frames[5][26][2] = 8'hac;
frames[5][26][3] = 8'hac;
frames[5][26][4] = 8'hac;
frames[5][26][5] = 8'hb1;
frames[5][26][6] = 8'hd1;
frames[5][26][7] = 8'hd1;
frames[5][26][8] = 8'hd1;
frames[5][26][9] = 8'hd1;
frames[5][26][10] = 8'hb1;
frames[5][26][11] = 8'hac;
frames[5][26][12] = 8'had;
frames[5][26][13] = 8'hb1;
frames[5][26][14] = 8'hb1;
frames[5][26][15] = 8'hb1;
frames[5][26][16] = 8'hb1;
frames[5][26][17] = 8'hb1;
frames[5][26][18] = 8'hd1;
frames[5][26][19] = 8'hd6;
frames[5][26][20] = 8'hd6;
frames[5][26][21] = 8'hd6;
frames[5][26][22] = 8'hd6;
frames[5][26][23] = 8'hd6;
frames[5][26][24] = 8'hd1;
frames[5][26][25] = 8'hd1;
frames[5][26][26] = 8'hd1;
frames[5][26][27] = 8'hb1;
frames[5][26][28] = 8'hb1;
frames[5][26][29] = 8'hb1;
frames[5][26][30] = 8'hb1;
frames[5][26][31] = 8'hb1;
frames[5][26][32] = 8'hb1;
frames[5][26][33] = 8'hb1;
frames[5][26][34] = 8'hb1;
frames[5][26][35] = 8'hb1;
frames[5][26][36] = 8'hb1;
frames[5][26][37] = 8'hb1;
frames[5][26][38] = 8'hb1;
frames[5][26][39] = 8'hb1;
frames[5][27][0] = 8'h8c;
frames[5][27][1] = 8'h8c;
frames[5][27][2] = 8'h8c;
frames[5][27][3] = 8'hac;
frames[5][27][4] = 8'hac;
frames[5][27][5] = 8'hb1;
frames[5][27][6] = 8'hb1;
frames[5][27][7] = 8'hb1;
frames[5][27][8] = 8'hd1;
frames[5][27][9] = 8'hd1;
frames[5][27][10] = 8'hb1;
frames[5][27][11] = 8'hb1;
frames[5][27][12] = 8'had;
frames[5][27][13] = 8'hb1;
frames[5][27][14] = 8'hb1;
frames[5][27][15] = 8'hb1;
frames[5][27][16] = 8'hac;
frames[5][27][17] = 8'hac;
frames[5][27][18] = 8'hb1;
frames[5][27][19] = 8'hd5;
frames[5][27][20] = 8'hd6;
frames[5][27][21] = 8'hd6;
frames[5][27][22] = 8'hda;
frames[5][27][23] = 8'hd6;
frames[5][27][24] = 8'hd1;
frames[5][27][25] = 8'hb1;
frames[5][27][26] = 8'hd1;
frames[5][27][27] = 8'hb1;
frames[5][27][28] = 8'hb1;
frames[5][27][29] = 8'hb1;
frames[5][27][30] = 8'hb1;
frames[5][27][31] = 8'hb1;
frames[5][27][32] = 8'hb1;
frames[5][27][33] = 8'hb1;
frames[5][27][34] = 8'hb1;
frames[5][27][35] = 8'hb1;
frames[5][27][36] = 8'hb1;
frames[5][27][37] = 8'hb1;
frames[5][27][38] = 8'hb1;
frames[5][27][39] = 8'hb1;
frames[5][28][0] = 8'h88;
frames[5][28][1] = 8'h8c;
frames[5][28][2] = 8'h8c;
frames[5][28][3] = 8'h8c;
frames[5][28][4] = 8'hac;
frames[5][28][5] = 8'had;
frames[5][28][6] = 8'hb1;
frames[5][28][7] = 8'hb1;
frames[5][28][8] = 8'hd1;
frames[5][28][9] = 8'hd1;
frames[5][28][10] = 8'hb1;
frames[5][28][11] = 8'hb1;
frames[5][28][12] = 8'hb1;
frames[5][28][13] = 8'hb1;
frames[5][28][14] = 8'hb1;
frames[5][28][15] = 8'hb1;
frames[5][28][16] = 8'hac;
frames[5][28][17] = 8'h8c;
frames[5][28][18] = 8'had;
frames[5][28][19] = 8'had;
frames[5][28][20] = 8'had;
frames[5][28][21] = 8'hb1;
frames[5][28][22] = 8'hd1;
frames[5][28][23] = 8'hd1;
frames[5][28][24] = 8'hb1;
frames[5][28][25] = 8'hb1;
frames[5][28][26] = 8'hb1;
frames[5][28][27] = 8'hb1;
frames[5][28][28] = 8'hb1;
frames[5][28][29] = 8'hb1;
frames[5][28][30] = 8'hb1;
frames[5][28][31] = 8'hb1;
frames[5][28][32] = 8'hb1;
frames[5][28][33] = 8'hb1;
frames[5][28][34] = 8'hb1;
frames[5][28][35] = 8'hb1;
frames[5][28][36] = 8'hb1;
frames[5][28][37] = 8'hb1;
frames[5][28][38] = 8'hb1;
frames[5][28][39] = 8'hb1;
frames[5][29][0] = 8'h88;
frames[5][29][1] = 8'h8c;
frames[5][29][2] = 8'h8c;
frames[5][29][3] = 8'h8c;
frames[5][29][4] = 8'hac;
frames[5][29][5] = 8'hac;
frames[5][29][6] = 8'hac;
frames[5][29][7] = 8'hb1;
frames[5][29][8] = 8'hd1;
frames[5][29][9] = 8'hd1;
frames[5][29][10] = 8'hb1;
frames[5][29][11] = 8'hb1;
frames[5][29][12] = 8'had;
frames[5][29][13] = 8'hb1;
frames[5][29][14] = 8'hb1;
frames[5][29][15] = 8'hb1;
frames[5][29][16] = 8'hac;
frames[5][29][17] = 8'h8c;
frames[5][29][18] = 8'h8c;
frames[5][29][19] = 8'h8c;
frames[5][29][20] = 8'h8c;
frames[5][29][21] = 8'h8c;
frames[5][29][22] = 8'had;
frames[5][29][23] = 8'hb1;
frames[5][29][24] = 8'hb1;
frames[5][29][25] = 8'hb1;
frames[5][29][26] = 8'hb1;
frames[5][29][27] = 8'hb1;
frames[5][29][28] = 8'hb1;
frames[5][29][29] = 8'hb1;
frames[5][29][30] = 8'hb1;
frames[5][29][31] = 8'hb1;
frames[5][29][32] = 8'hb1;
frames[5][29][33] = 8'hb1;
frames[5][29][34] = 8'hb1;
frames[5][29][35] = 8'hb1;
frames[5][29][36] = 8'hb1;
frames[5][29][37] = 8'hb1;
frames[5][29][38] = 8'hb1;
frames[5][29][39] = 8'hb1;
frames[6][0][0] = 8'hb1;
frames[6][0][1] = 8'hb1;
frames[6][0][2] = 8'hb1;
frames[6][0][3] = 8'hd1;
frames[6][0][4] = 8'hd1;
frames[6][0][5] = 8'hd1;
frames[6][0][6] = 8'hd1;
frames[6][0][7] = 8'hd5;
frames[6][0][8] = 8'hd1;
frames[6][0][9] = 8'hd1;
frames[6][0][10] = 8'hd1;
frames[6][0][11] = 8'hd5;
frames[6][0][12] = 8'hd5;
frames[6][0][13] = 8'hd5;
frames[6][0][14] = 8'hd5;
frames[6][0][15] = 8'hd5;
frames[6][0][16] = 8'hd5;
frames[6][0][17] = 8'hd1;
frames[6][0][18] = 8'hd1;
frames[6][0][19] = 8'hd1;
frames[6][0][20] = 8'hd1;
frames[6][0][21] = 8'hd1;
frames[6][0][22] = 8'hd5;
frames[6][0][23] = 8'hd5;
frames[6][0][24] = 8'hd5;
frames[6][0][25] = 8'hd5;
frames[6][0][26] = 8'hd5;
frames[6][0][27] = 8'hd1;
frames[6][0][28] = 8'hd1;
frames[6][0][29] = 8'hd1;
frames[6][0][30] = 8'hd1;
frames[6][0][31] = 8'hd1;
frames[6][0][32] = 8'hd1;
frames[6][0][33] = 8'hd5;
frames[6][0][34] = 8'hd1;
frames[6][0][35] = 8'hd1;
frames[6][0][36] = 8'hd1;
frames[6][0][37] = 8'hd1;
frames[6][0][38] = 8'hb1;
frames[6][0][39] = 8'had;
frames[6][1][0] = 8'hb1;
frames[6][1][1] = 8'hb1;
frames[6][1][2] = 8'hb1;
frames[6][1][3] = 8'hd1;
frames[6][1][4] = 8'hd1;
frames[6][1][5] = 8'hd1;
frames[6][1][6] = 8'hd1;
frames[6][1][7] = 8'hd1;
frames[6][1][8] = 8'hd1;
frames[6][1][9] = 8'hd1;
frames[6][1][10] = 8'hd1;
frames[6][1][11] = 8'hd5;
frames[6][1][12] = 8'hd5;
frames[6][1][13] = 8'hd5;
frames[6][1][14] = 8'hd5;
frames[6][1][15] = 8'hd5;
frames[6][1][16] = 8'hd5;
frames[6][1][17] = 8'hd1;
frames[6][1][18] = 8'hd1;
frames[6][1][19] = 8'hd1;
frames[6][1][20] = 8'hd1;
frames[6][1][21] = 8'hd1;
frames[6][1][22] = 8'hd5;
frames[6][1][23] = 8'hd5;
frames[6][1][24] = 8'hd5;
frames[6][1][25] = 8'hd5;
frames[6][1][26] = 8'hd5;
frames[6][1][27] = 8'hd1;
frames[6][1][28] = 8'hd1;
frames[6][1][29] = 8'hd1;
frames[6][1][30] = 8'hd1;
frames[6][1][31] = 8'hd1;
frames[6][1][32] = 8'hd1;
frames[6][1][33] = 8'hd5;
frames[6][1][34] = 8'hd1;
frames[6][1][35] = 8'hd1;
frames[6][1][36] = 8'hd1;
frames[6][1][37] = 8'hd1;
frames[6][1][38] = 8'hb1;
frames[6][1][39] = 8'had;
frames[6][2][0] = 8'hb1;
frames[6][2][1] = 8'hb1;
frames[6][2][2] = 8'hd1;
frames[6][2][3] = 8'hd1;
frames[6][2][4] = 8'hd1;
frames[6][2][5] = 8'hd1;
frames[6][2][6] = 8'hd5;
frames[6][2][7] = 8'hd5;
frames[6][2][8] = 8'hd5;
frames[6][2][9] = 8'hd5;
frames[6][2][10] = 8'hd5;
frames[6][2][11] = 8'hd5;
frames[6][2][12] = 8'hf5;
frames[6][2][13] = 8'hd5;
frames[6][2][14] = 8'hd5;
frames[6][2][15] = 8'hd5;
frames[6][2][16] = 8'hd1;
frames[6][2][17] = 8'hd1;
frames[6][2][18] = 8'hd1;
frames[6][2][19] = 8'hd1;
frames[6][2][20] = 8'hd1;
frames[6][2][21] = 8'hd1;
frames[6][2][22] = 8'hd5;
frames[6][2][23] = 8'hd5;
frames[6][2][24] = 8'hd5;
frames[6][2][25] = 8'hd5;
frames[6][2][26] = 8'hd5;
frames[6][2][27] = 8'hd1;
frames[6][2][28] = 8'hd1;
frames[6][2][29] = 8'hd1;
frames[6][2][30] = 8'hd1;
frames[6][2][31] = 8'hd1;
frames[6][2][32] = 8'hd1;
frames[6][2][33] = 8'hd1;
frames[6][2][34] = 8'hd1;
frames[6][2][35] = 8'hd1;
frames[6][2][36] = 8'hd1;
frames[6][2][37] = 8'hd1;
frames[6][2][38] = 8'hb1;
frames[6][2][39] = 8'hac;
frames[6][3][0] = 8'hb1;
frames[6][3][1] = 8'hb1;
frames[6][3][2] = 8'hd1;
frames[6][3][3] = 8'hd1;
frames[6][3][4] = 8'hd1;
frames[6][3][5] = 8'hd1;
frames[6][3][6] = 8'hd6;
frames[6][3][7] = 8'hd6;
frames[6][3][8] = 8'hd6;
frames[6][3][9] = 8'hd6;
frames[6][3][10] = 8'hd6;
frames[6][3][11] = 8'hd6;
frames[6][3][12] = 8'hf6;
frames[6][3][13] = 8'hd5;
frames[6][3][14] = 8'hd5;
frames[6][3][15] = 8'hd5;
frames[6][3][16] = 8'hd1;
frames[6][3][17] = 8'hd1;
frames[6][3][18] = 8'hd1;
frames[6][3][19] = 8'hd1;
frames[6][3][20] = 8'hd1;
frames[6][3][21] = 8'hd1;
frames[6][3][22] = 8'hd5;
frames[6][3][23] = 8'hd5;
frames[6][3][24] = 8'hd5;
frames[6][3][25] = 8'hd5;
frames[6][3][26] = 8'hd5;
frames[6][3][27] = 8'hd1;
frames[6][3][28] = 8'hd1;
frames[6][3][29] = 8'hd1;
frames[6][3][30] = 8'hd1;
frames[6][3][31] = 8'hd1;
frames[6][3][32] = 8'hd1;
frames[6][3][33] = 8'hd5;
frames[6][3][34] = 8'hd1;
frames[6][3][35] = 8'hd1;
frames[6][3][36] = 8'hd1;
frames[6][3][37] = 8'hd1;
frames[6][3][38] = 8'hb1;
frames[6][3][39] = 8'hac;
frames[6][4][0] = 8'hb1;
frames[6][4][1] = 8'hb1;
frames[6][4][2] = 8'hd1;
frames[6][4][3] = 8'hd1;
frames[6][4][4] = 8'hd1;
frames[6][4][5] = 8'hd1;
frames[6][4][6] = 8'hd1;
frames[6][4][7] = 8'hd5;
frames[6][4][8] = 8'hd5;
frames[6][4][9] = 8'hd1;
frames[6][4][10] = 8'hd5;
frames[6][4][11] = 8'hd5;
frames[6][4][12] = 8'hd5;
frames[6][4][13] = 8'hd5;
frames[6][4][14] = 8'hd5;
frames[6][4][15] = 8'hd5;
frames[6][4][16] = 8'hd1;
frames[6][4][17] = 8'hd1;
frames[6][4][18] = 8'hd1;
frames[6][4][19] = 8'hd1;
frames[6][4][20] = 8'hd1;
frames[6][4][21] = 8'hd1;
frames[6][4][22] = 8'hd5;
frames[6][4][23] = 8'hd1;
frames[6][4][24] = 8'hd1;
frames[6][4][25] = 8'hd1;
frames[6][4][26] = 8'hd1;
frames[6][4][27] = 8'hd1;
frames[6][4][28] = 8'hd1;
frames[6][4][29] = 8'hd1;
frames[6][4][30] = 8'hd1;
frames[6][4][31] = 8'hd1;
frames[6][4][32] = 8'hd1;
frames[6][4][33] = 8'hd5;
frames[6][4][34] = 8'hd5;
frames[6][4][35] = 8'hd1;
frames[6][4][36] = 8'hd1;
frames[6][4][37] = 8'hd1;
frames[6][4][38] = 8'hd1;
frames[6][4][39] = 8'hb0;
frames[6][5][0] = 8'hb1;
frames[6][5][1] = 8'hb1;
frames[6][5][2] = 8'hb1;
frames[6][5][3] = 8'hd1;
frames[6][5][4] = 8'hd1;
frames[6][5][5] = 8'hd1;
frames[6][5][6] = 8'hd1;
frames[6][5][7] = 8'hd1;
frames[6][5][8] = 8'hd1;
frames[6][5][9] = 8'hb1;
frames[6][5][10] = 8'hb1;
frames[6][5][11] = 8'hd1;
frames[6][5][12] = 8'hd5;
frames[6][5][13] = 8'hd5;
frames[6][5][14] = 8'hd1;
frames[6][5][15] = 8'hd5;
frames[6][5][16] = 8'hd1;
frames[6][5][17] = 8'hd1;
frames[6][5][18] = 8'hd1;
frames[6][5][19] = 8'hd1;
frames[6][5][20] = 8'hd1;
frames[6][5][21] = 8'hd1;
frames[6][5][22] = 8'hd1;
frames[6][5][23] = 8'hd1;
frames[6][5][24] = 8'hd1;
frames[6][5][25] = 8'hd1;
frames[6][5][26] = 8'hd1;
frames[6][5][27] = 8'hd1;
frames[6][5][28] = 8'hd1;
frames[6][5][29] = 8'hd1;
frames[6][5][30] = 8'hd5;
frames[6][5][31] = 8'hd5;
frames[6][5][32] = 8'hd5;
frames[6][5][33] = 8'hd5;
frames[6][5][34] = 8'hd5;
frames[6][5][35] = 8'hd5;
frames[6][5][36] = 8'hd1;
frames[6][5][37] = 8'hd1;
frames[6][5][38] = 8'hd1;
frames[6][5][39] = 8'hac;
frames[6][6][0] = 8'hb1;
frames[6][6][1] = 8'hb1;
frames[6][6][2] = 8'hb1;
frames[6][6][3] = 8'hd1;
frames[6][6][4] = 8'hd1;
frames[6][6][5] = 8'hd1;
frames[6][6][6] = 8'hd1;
frames[6][6][7] = 8'hd5;
frames[6][6][8] = 8'hd1;
frames[6][6][9] = 8'hb1;
frames[6][6][10] = 8'hd1;
frames[6][6][11] = 8'hfa;
frames[6][6][12] = 8'hda;
frames[6][6][13] = 8'hda;
frames[6][6][14] = 8'hfa;
frames[6][6][15] = 8'hd5;
frames[6][6][16] = 8'hb1;
frames[6][6][17] = 8'hd6;
frames[6][6][18] = 8'hb1;
frames[6][6][19] = 8'h91;
frames[6][6][20] = 8'h8d;
frames[6][6][21] = 8'hb6;
frames[6][6][22] = 8'hb6;
frames[6][6][23] = 8'h96;
frames[6][6][24] = 8'hb6;
frames[6][6][25] = 8'h96;
frames[6][6][26] = 8'h91;
frames[6][6][27] = 8'h6d;
frames[6][6][28] = 8'h68;
frames[6][6][29] = 8'hd1;
frames[6][6][30] = 8'hd5;
frames[6][6][31] = 8'hd6;
frames[6][6][32] = 8'hd6;
frames[6][6][33] = 8'hd6;
frames[6][6][34] = 8'hd6;
frames[6][6][35] = 8'hd5;
frames[6][6][36] = 8'hd1;
frames[6][6][37] = 8'hd1;
frames[6][6][38] = 8'hd1;
frames[6][6][39] = 8'hac;
frames[6][7][0] = 8'hb1;
frames[6][7][1] = 8'hb1;
frames[6][7][2] = 8'hd1;
frames[6][7][3] = 8'hd1;
frames[6][7][4] = 8'hd1;
frames[6][7][5] = 8'hd1;
frames[6][7][6] = 8'hd1;
frames[6][7][7] = 8'hd1;
frames[6][7][8] = 8'hd1;
frames[6][7][9] = 8'hd1;
frames[6][7][10] = 8'hd6;
frames[6][7][11] = 8'hfe;
frames[6][7][12] = 8'hfe;
frames[6][7][13] = 8'hfe;
frames[6][7][14] = 8'hfe;
frames[6][7][15] = 8'hd6;
frames[6][7][16] = 8'hb1;
frames[6][7][17] = 8'hb1;
frames[6][7][18] = 8'h8d;
frames[6][7][19] = 8'h69;
frames[6][7][20] = 8'h96;
frames[6][7][21] = 8'h96;
frames[6][7][22] = 8'hb6;
frames[6][7][23] = 8'hda;
frames[6][7][24] = 8'hda;
frames[6][7][25] = 8'hb6;
frames[6][7][26] = 8'h92;
frames[6][7][27] = 8'h49;
frames[6][7][28] = 8'h20;
frames[6][7][29] = 8'hb1;
frames[6][7][30] = 8'hd5;
frames[6][7][31] = 8'hd5;
frames[6][7][32] = 8'hd5;
frames[6][7][33] = 8'hd5;
frames[6][7][34] = 8'hd5;
frames[6][7][35] = 8'hd5;
frames[6][7][36] = 8'hd1;
frames[6][7][37] = 8'hd1;
frames[6][7][38] = 8'hd1;
frames[6][7][39] = 8'had;
frames[6][8][0] = 8'hac;
frames[6][8][1] = 8'hb1;
frames[6][8][2] = 8'hb1;
frames[6][8][3] = 8'hb1;
frames[6][8][4] = 8'hb1;
frames[6][8][5] = 8'hb1;
frames[6][8][6] = 8'hd1;
frames[6][8][7] = 8'hd1;
frames[6][8][8] = 8'hd1;
frames[6][8][9] = 8'hd5;
frames[6][8][10] = 8'hfa;
frames[6][8][11] = 8'hfa;
frames[6][8][12] = 8'hfa;
frames[6][8][13] = 8'hfa;
frames[6][8][14] = 8'hfa;
frames[6][8][15] = 8'hfa;
frames[6][8][16] = 8'hb1;
frames[6][8][17] = 8'h91;
frames[6][8][18] = 8'h6d;
frames[6][8][19] = 8'hb6;
frames[6][8][20] = 8'hb6;
frames[6][8][21] = 8'hda;
frames[6][8][22] = 8'hfa;
frames[6][8][23] = 8'hfa;
frames[6][8][24] = 8'hfa;
frames[6][8][25] = 8'hfa;
frames[6][8][26] = 8'hba;
frames[6][8][27] = 8'h92;
frames[6][8][28] = 8'h44;
frames[6][8][29] = 8'hb1;
frames[6][8][30] = 8'hd1;
frames[6][8][31] = 8'hd5;
frames[6][8][32] = 8'hd1;
frames[6][8][33] = 8'hd5;
frames[6][8][34] = 8'hd5;
frames[6][8][35] = 8'hd5;
frames[6][8][36] = 8'hd1;
frames[6][8][37] = 8'hd1;
frames[6][8][38] = 8'hd1;
frames[6][8][39] = 8'had;
frames[6][9][0] = 8'hac;
frames[6][9][1] = 8'hb1;
frames[6][9][2] = 8'hb1;
frames[6][9][3] = 8'hb1;
frames[6][9][4] = 8'hb1;
frames[6][9][5] = 8'hb1;
frames[6][9][6] = 8'hd1;
frames[6][9][7] = 8'hd1;
frames[6][9][8] = 8'hb1;
frames[6][9][9] = 8'hb1;
frames[6][9][10] = 8'hd6;
frames[6][9][11] = 8'hfa;
frames[6][9][12] = 8'hfa;
frames[6][9][13] = 8'hfa;
frames[6][9][14] = 8'hfa;
frames[6][9][15] = 8'hfa;
frames[6][9][16] = 8'hb6;
frames[6][9][17] = 8'h91;
frames[6][9][18] = 8'h92;
frames[6][9][19] = 8'hda;
frames[6][9][20] = 8'hfa;
frames[6][9][21] = 8'hfa;
frames[6][9][22] = 8'hfa;
frames[6][9][23] = 8'hfa;
frames[6][9][24] = 8'hfa;
frames[6][9][25] = 8'hfa;
frames[6][9][26] = 8'hff;
frames[6][9][27] = 8'hda;
frames[6][9][28] = 8'h91;
frames[6][9][29] = 8'hb1;
frames[6][9][30] = 8'hf5;
frames[6][9][31] = 8'hd1;
frames[6][9][32] = 8'hd1;
frames[6][9][33] = 8'hd1;
frames[6][9][34] = 8'hd5;
frames[6][9][35] = 8'hd5;
frames[6][9][36] = 8'hd1;
frames[6][9][37] = 8'hd1;
frames[6][9][38] = 8'hd1;
frames[6][9][39] = 8'hb1;
frames[6][10][0] = 8'hac;
frames[6][10][1] = 8'hb1;
frames[6][10][2] = 8'hb1;
frames[6][10][3] = 8'hb1;
frames[6][10][4] = 8'hb1;
frames[6][10][5] = 8'hb1;
frames[6][10][6] = 8'hd1;
frames[6][10][7] = 8'hd1;
frames[6][10][8] = 8'hb1;
frames[6][10][9] = 8'had;
frames[6][10][10] = 8'hd6;
frames[6][10][11] = 8'hfa;
frames[6][10][12] = 8'hfa;
frames[6][10][13] = 8'hfa;
frames[6][10][14] = 8'hfa;
frames[6][10][15] = 8'hfa;
frames[6][10][16] = 8'hb6;
frames[6][10][17] = 8'h91;
frames[6][10][18] = 8'hd6;
frames[6][10][19] = 8'hff;
frames[6][10][20] = 8'hfa;
frames[6][10][21] = 8'hfa;
frames[6][10][22] = 8'hfa;
frames[6][10][23] = 8'hfa;
frames[6][10][24] = 8'hfa;
frames[6][10][25] = 8'hfa;
frames[6][10][26] = 8'hfb;
frames[6][10][27] = 8'hfb;
frames[6][10][28] = 8'hda;
frames[6][10][29] = 8'hb6;
frames[6][10][30] = 8'hd1;
frames[6][10][31] = 8'hd1;
frames[6][10][32] = 8'hd1;
frames[6][10][33] = 8'hd1;
frames[6][10][34] = 8'hd5;
frames[6][10][35] = 8'hd5;
frames[6][10][36] = 8'hd1;
frames[6][10][37] = 8'hb1;
frames[6][10][38] = 8'hd1;
frames[6][10][39] = 8'hb1;
frames[6][11][0] = 8'hac;
frames[6][11][1] = 8'hac;
frames[6][11][2] = 8'hb1;
frames[6][11][3] = 8'hb1;
frames[6][11][4] = 8'hb1;
frames[6][11][5] = 8'hd1;
frames[6][11][6] = 8'hd1;
frames[6][11][7] = 8'hd1;
frames[6][11][8] = 8'hb1;
frames[6][11][9] = 8'had;
frames[6][11][10] = 8'hd5;
frames[6][11][11] = 8'hda;
frames[6][11][12] = 8'hda;
frames[6][11][13] = 8'hfa;
frames[6][11][14] = 8'hfa;
frames[6][11][15] = 8'hfa;
frames[6][11][16] = 8'hb2;
frames[6][11][17] = 8'hb2;
frames[6][11][18] = 8'hfa;
frames[6][11][19] = 8'hff;
frames[6][11][20] = 8'hfa;
frames[6][11][21] = 8'hfa;
frames[6][11][22] = 8'hfa;
frames[6][11][23] = 8'hfa;
frames[6][11][24] = 8'hfa;
frames[6][11][25] = 8'hfa;
frames[6][11][26] = 8'hfa;
frames[6][11][27] = 8'hfa;
frames[6][11][28] = 8'hda;
frames[6][11][29] = 8'hb6;
frames[6][11][30] = 8'hd1;
frames[6][11][31] = 8'hd1;
frames[6][11][32] = 8'hd1;
frames[6][11][33] = 8'hd1;
frames[6][11][34] = 8'hd5;
frames[6][11][35] = 8'hd5;
frames[6][11][36] = 8'hd1;
frames[6][11][37] = 8'hb1;
frames[6][11][38] = 8'hb1;
frames[6][11][39] = 8'hb1;
frames[6][12][0] = 8'hac;
frames[6][12][1] = 8'had;
frames[6][12][2] = 8'hb1;
frames[6][12][3] = 8'hb1;
frames[6][12][4] = 8'hb1;
frames[6][12][5] = 8'hb1;
frames[6][12][6] = 8'hb1;
frames[6][12][7] = 8'hb1;
frames[6][12][8] = 8'hb1;
frames[6][12][9] = 8'had;
frames[6][12][10] = 8'hb1;
frames[6][12][11] = 8'hd6;
frames[6][12][12] = 8'hfa;
frames[6][12][13] = 8'hfa;
frames[6][12][14] = 8'hfa;
frames[6][12][15] = 8'hd6;
frames[6][12][16] = 8'hb1;
frames[6][12][17] = 8'hb6;
frames[6][12][18] = 8'hfa;
frames[6][12][19] = 8'hfb;
frames[6][12][20] = 8'hfb;
frames[6][12][21] = 8'hfa;
frames[6][12][22] = 8'hfa;
frames[6][12][23] = 8'hfa;
frames[6][12][24] = 8'hfa;
frames[6][12][25] = 8'hfa;
frames[6][12][26] = 8'hfa;
frames[6][12][27] = 8'hfa;
frames[6][12][28] = 8'hfa;
frames[6][12][29] = 8'hb6;
frames[6][12][30] = 8'hd1;
frames[6][12][31] = 8'hd1;
frames[6][12][32] = 8'hd1;
frames[6][12][33] = 8'hd1;
frames[6][12][34] = 8'hd5;
frames[6][12][35] = 8'hd5;
frames[6][12][36] = 8'hd1;
frames[6][12][37] = 8'hb1;
frames[6][12][38] = 8'hb1;
frames[6][12][39] = 8'hb1;
frames[6][13][0] = 8'hac;
frames[6][13][1] = 8'hac;
frames[6][13][2] = 8'hb1;
frames[6][13][3] = 8'hb0;
frames[6][13][4] = 8'hb1;
frames[6][13][5] = 8'hb1;
frames[6][13][6] = 8'hb1;
frames[6][13][7] = 8'hb1;
frames[6][13][8] = 8'had;
frames[6][13][9] = 8'hac;
frames[6][13][10] = 8'h8d;
frames[6][13][11] = 8'hb1;
frames[6][13][12] = 8'hd6;
frames[6][13][13] = 8'hfa;
frames[6][13][14] = 8'hda;
frames[6][13][15] = 8'hb1;
frames[6][13][16] = 8'h91;
frames[6][13][17] = 8'hb6;
frames[6][13][18] = 8'hfa;
frames[6][13][19] = 8'hff;
frames[6][13][20] = 8'hfb;
frames[6][13][21] = 8'hfb;
frames[6][13][22] = 8'hfa;
frames[6][13][23] = 8'hfa;
frames[6][13][24] = 8'hfa;
frames[6][13][25] = 8'hfa;
frames[6][13][26] = 8'hfa;
frames[6][13][27] = 8'hfa;
frames[6][13][28] = 8'hfa;
frames[6][13][29] = 8'hd6;
frames[6][13][30] = 8'hd1;
frames[6][13][31] = 8'hd1;
frames[6][13][32] = 8'hd1;
frames[6][13][33] = 8'hd1;
frames[6][13][34] = 8'hd5;
frames[6][13][35] = 8'hd5;
frames[6][13][36] = 8'hd1;
frames[6][13][37] = 8'hb1;
frames[6][13][38] = 8'hb1;
frames[6][13][39] = 8'hb1;
frames[6][14][0] = 8'hac;
frames[6][14][1] = 8'hac;
frames[6][14][2] = 8'hb1;
frames[6][14][3] = 8'hb1;
frames[6][14][4] = 8'hb1;
frames[6][14][5] = 8'hb1;
frames[6][14][6] = 8'hb1;
frames[6][14][7] = 8'hac;
frames[6][14][8] = 8'had;
frames[6][14][9] = 8'hac;
frames[6][14][10] = 8'h8d;
frames[6][14][11] = 8'h91;
frames[6][14][12] = 8'hb1;
frames[6][14][13] = 8'hb5;
frames[6][14][14] = 8'h91;
frames[6][14][15] = 8'hb1;
frames[6][14][16] = 8'h91;
frames[6][14][17] = 8'h91;
frames[6][14][18] = 8'hfa;
frames[6][14][19] = 8'hff;
frames[6][14][20] = 8'hff;
frames[6][14][21] = 8'hfa;
frames[6][14][22] = 8'hfa;
frames[6][14][23] = 8'hfa;
frames[6][14][24] = 8'hfa;
frames[6][14][25] = 8'hfa;
frames[6][14][26] = 8'hfa;
frames[6][14][27] = 8'hfa;
frames[6][14][28] = 8'hfa;
frames[6][14][29] = 8'hb6;
frames[6][14][30] = 8'hd1;
frames[6][14][31] = 8'hd1;
frames[6][14][32] = 8'hd1;
frames[6][14][33] = 8'hd1;
frames[6][14][34] = 8'hd1;
frames[6][14][35] = 8'hd5;
frames[6][14][36] = 8'hd1;
frames[6][14][37] = 8'hb1;
frames[6][14][38] = 8'hb1;
frames[6][14][39] = 8'hb1;
frames[6][15][0] = 8'hac;
frames[6][15][1] = 8'hac;
frames[6][15][2] = 8'hac;
frames[6][15][3] = 8'hac;
frames[6][15][4] = 8'hac;
frames[6][15][5] = 8'hb1;
frames[6][15][6] = 8'hb1;
frames[6][15][7] = 8'hac;
frames[6][15][8] = 8'hac;
frames[6][15][9] = 8'hac;
frames[6][15][10] = 8'h8d;
frames[6][15][11] = 8'h89;
frames[6][15][12] = 8'h89;
frames[6][15][13] = 8'h8d;
frames[6][15][14] = 8'h91;
frames[6][15][15] = 8'h91;
frames[6][15][16] = 8'h8d;
frames[6][15][17] = 8'h8d;
frames[6][15][18] = 8'hfa;
frames[6][15][19] = 8'hff;
frames[6][15][20] = 8'hfb;
frames[6][15][21] = 8'hfb;
frames[6][15][22] = 8'hfa;
frames[6][15][23] = 8'hfa;
frames[6][15][24] = 8'hfa;
frames[6][15][25] = 8'hfa;
frames[6][15][26] = 8'hfa;
frames[6][15][27] = 8'hfa;
frames[6][15][28] = 8'hda;
frames[6][15][29] = 8'hb6;
frames[6][15][30] = 8'hd1;
frames[6][15][31] = 8'hd1;
frames[6][15][32] = 8'hd1;
frames[6][15][33] = 8'hd1;
frames[6][15][34] = 8'hd1;
frames[6][15][35] = 8'hd5;
frames[6][15][36] = 8'hd1;
frames[6][15][37] = 8'hb1;
frames[6][15][38] = 8'hb1;
frames[6][15][39] = 8'hb1;
frames[6][16][0] = 8'hac;
frames[6][16][1] = 8'hac;
frames[6][16][2] = 8'hac;
frames[6][16][3] = 8'hac;
frames[6][16][4] = 8'hac;
frames[6][16][5] = 8'hb1;
frames[6][16][6] = 8'hb1;
frames[6][16][7] = 8'hac;
frames[6][16][8] = 8'hac;
frames[6][16][9] = 8'h8c;
frames[6][16][10] = 8'had;
frames[6][16][11] = 8'h64;
frames[6][16][12] = 8'h60;
frames[6][16][13] = 8'h84;
frames[6][16][14] = 8'h8d;
frames[6][16][15] = 8'hb1;
frames[6][16][16] = 8'h91;
frames[6][16][17] = 8'h8d;
frames[6][16][18] = 8'hd6;
frames[6][16][19] = 8'hff;
frames[6][16][20] = 8'hfa;
frames[6][16][21] = 8'hfa;
frames[6][16][22] = 8'hfa;
frames[6][16][23] = 8'hfa;
frames[6][16][24] = 8'hfa;
frames[6][16][25] = 8'hfa;
frames[6][16][26] = 8'hfa;
frames[6][16][27] = 8'hfa;
frames[6][16][28] = 8'hda;
frames[6][16][29] = 8'h91;
frames[6][16][30] = 8'hb1;
frames[6][16][31] = 8'hd1;
frames[6][16][32] = 8'hd1;
frames[6][16][33] = 8'hd1;
frames[6][16][34] = 8'hd1;
frames[6][16][35] = 8'hd5;
frames[6][16][36] = 8'hd1;
frames[6][16][37] = 8'hb1;
frames[6][16][38] = 8'hb1;
frames[6][16][39] = 8'hb1;
frames[6][17][0] = 8'hac;
frames[6][17][1] = 8'hac;
frames[6][17][2] = 8'hac;
frames[6][17][3] = 8'hac;
frames[6][17][4] = 8'hac;
frames[6][17][5] = 8'hb1;
frames[6][17][6] = 8'hb1;
frames[6][17][7] = 8'hac;
frames[6][17][8] = 8'hac;
frames[6][17][9] = 8'h8c;
frames[6][17][10] = 8'h84;
frames[6][17][11] = 8'h60;
frames[6][17][12] = 8'h60;
frames[6][17][13] = 8'h60;
frames[6][17][14] = 8'h69;
frames[6][17][15] = 8'h8d;
frames[6][17][16] = 8'h91;
frames[6][17][17] = 8'h8d;
frames[6][17][18] = 8'hb1;
frames[6][17][19] = 8'hfb;
frames[6][17][20] = 8'hfb;
frames[6][17][21] = 8'hfa;
frames[6][17][22] = 8'hfa;
frames[6][17][23] = 8'hfa;
frames[6][17][24] = 8'hfa;
frames[6][17][25] = 8'hfa;
frames[6][17][26] = 8'hfa;
frames[6][17][27] = 8'hfa;
frames[6][17][28] = 8'hb6;
frames[6][17][29] = 8'h6d;
frames[6][17][30] = 8'hb1;
frames[6][17][31] = 8'hd1;
frames[6][17][32] = 8'hd1;
frames[6][17][33] = 8'hd1;
frames[6][17][34] = 8'hd1;
frames[6][17][35] = 8'hd1;
frames[6][17][36] = 8'hd1;
frames[6][17][37] = 8'hb1;
frames[6][17][38] = 8'hb1;
frames[6][17][39] = 8'hb1;
frames[6][18][0] = 8'hac;
frames[6][18][1] = 8'hac;
frames[6][18][2] = 8'hac;
frames[6][18][3] = 8'hac;
frames[6][18][4] = 8'hb0;
frames[6][18][5] = 8'hd1;
frames[6][18][6] = 8'hd1;
frames[6][18][7] = 8'hb1;
frames[6][18][8] = 8'had;
frames[6][18][9] = 8'h8c;
frames[6][18][10] = 8'h64;
frames[6][18][11] = 8'h60;
frames[6][18][12] = 8'h60;
frames[6][18][13] = 8'h60;
frames[6][18][14] = 8'h68;
frames[6][18][15] = 8'h8d;
frames[6][18][16] = 8'h8d;
frames[6][18][17] = 8'h8d;
frames[6][18][18] = 8'h6d;
frames[6][18][19] = 8'hd6;
frames[6][18][20] = 8'hfa;
frames[6][18][21] = 8'hfa;
frames[6][18][22] = 8'hfa;
frames[6][18][23] = 8'hfa;
frames[6][18][24] = 8'hfa;
frames[6][18][25] = 8'hfa;
frames[6][18][26] = 8'hda;
frames[6][18][27] = 8'hda;
frames[6][18][28] = 8'hb6;
frames[6][18][29] = 8'h48;
frames[6][18][30] = 8'hb1;
frames[6][18][31] = 8'hd1;
frames[6][18][32] = 8'hd1;
frames[6][18][33] = 8'hd1;
frames[6][18][34] = 8'hd1;
frames[6][18][35] = 8'hd1;
frames[6][18][36] = 8'hd1;
frames[6][18][37] = 8'hb1;
frames[6][18][38] = 8'hb1;
frames[6][18][39] = 8'hb1;
frames[6][19][0] = 8'hac;
frames[6][19][1] = 8'hac;
frames[6][19][2] = 8'hac;
frames[6][19][3] = 8'hac;
frames[6][19][4] = 8'hb0;
frames[6][19][5] = 8'hd1;
frames[6][19][6] = 8'hd1;
frames[6][19][7] = 8'hd1;
frames[6][19][8] = 8'hac;
frames[6][19][9] = 8'h8c;
frames[6][19][10] = 8'h84;
frames[6][19][11] = 8'h40;
frames[6][19][12] = 8'h60;
frames[6][19][13] = 8'h60;
frames[6][19][14] = 8'h68;
frames[6][19][15] = 8'h8d;
frames[6][19][16] = 8'h8d;
frames[6][19][17] = 8'h69;
frames[6][19][18] = 8'h68;
frames[6][19][19] = 8'h8d;
frames[6][19][20] = 8'hda;
frames[6][19][21] = 8'hdb;
frames[6][19][22] = 8'hfa;
frames[6][19][23] = 8'hda;
frames[6][19][24] = 8'hda;
frames[6][19][25] = 8'hda;
frames[6][19][26] = 8'hda;
frames[6][19][27] = 8'hb6;
frames[6][19][28] = 8'h8d;
frames[6][19][29] = 8'h44;
frames[6][19][30] = 8'hb1;
frames[6][19][31] = 8'hb1;
frames[6][19][32] = 8'hd1;
frames[6][19][33] = 8'hd1;
frames[6][19][34] = 8'hd1;
frames[6][19][35] = 8'hd1;
frames[6][19][36] = 8'hd1;
frames[6][19][37] = 8'hb1;
frames[6][19][38] = 8'hb1;
frames[6][19][39] = 8'hb1;
frames[6][20][0] = 8'hac;
frames[6][20][1] = 8'hac;
frames[6][20][2] = 8'hac;
frames[6][20][3] = 8'hac;
frames[6][20][4] = 8'hac;
frames[6][20][5] = 8'hb1;
frames[6][20][6] = 8'hd1;
frames[6][20][7] = 8'hb1;
frames[6][20][8] = 8'hac;
frames[6][20][9] = 8'had;
frames[6][20][10] = 8'h89;
frames[6][20][11] = 8'h64;
frames[6][20][12] = 8'h64;
frames[6][20][13] = 8'h88;
frames[6][20][14] = 8'h69;
frames[6][20][15] = 8'h8d;
frames[6][20][16] = 8'ha9;
frames[6][20][17] = 8'h88;
frames[6][20][18] = 8'ha8;
frames[6][20][19] = 8'ha4;
frames[6][20][20] = 8'h92;
frames[6][20][21] = 8'hba;
frames[6][20][22] = 8'hb6;
frames[6][20][23] = 8'h96;
frames[6][20][24] = 8'hb6;
frames[6][20][25] = 8'hba;
frames[6][20][26] = 8'hb6;
frames[6][20][27] = 8'hb6;
frames[6][20][28] = 8'h8d;
frames[6][20][29] = 8'h44;
frames[6][20][30] = 8'hb1;
frames[6][20][31] = 8'hb1;
frames[6][20][32] = 8'hd1;
frames[6][20][33] = 8'hd1;
frames[6][20][34] = 8'hd1;
frames[6][20][35] = 8'hd1;
frames[6][20][36] = 8'hb1;
frames[6][20][37] = 8'hb1;
frames[6][20][38] = 8'hb1;
frames[6][20][39] = 8'hb1;
frames[6][21][0] = 8'hac;
frames[6][21][1] = 8'hac;
frames[6][21][2] = 8'hb1;
frames[6][21][3] = 8'hd1;
frames[6][21][4] = 8'hd1;
frames[6][21][5] = 8'hd1;
frames[6][21][6] = 8'hd5;
frames[6][21][7] = 8'hd5;
frames[6][21][8] = 8'hb1;
frames[6][21][9] = 8'hb1;
frames[6][21][10] = 8'h8d;
frames[6][21][11] = 8'h8d;
frames[6][21][12] = 8'h91;
frames[6][21][13] = 8'h8d;
frames[6][21][14] = 8'h8d;
frames[6][21][15] = 8'h8d;
frames[6][21][16] = 8'ha8;
frames[6][21][17] = 8'h64;
frames[6][21][18] = 8'ha8;
frames[6][21][19] = 8'ha4;
frames[6][21][20] = 8'h8d;
frames[6][21][21] = 8'hb1;
frames[6][21][22] = 8'hb6;
frames[6][21][23] = 8'hb6;
frames[6][21][24] = 8'hb6;
frames[6][21][25] = 8'hb6;
frames[6][21][26] = 8'hb2;
frames[6][21][27] = 8'hb2;
frames[6][21][28] = 8'h91;
frames[6][21][29] = 8'h44;
frames[6][21][30] = 8'had;
frames[6][21][31] = 8'hb1;
frames[6][21][32] = 8'hd1;
frames[6][21][33] = 8'hd1;
frames[6][21][34] = 8'hb1;
frames[6][21][35] = 8'hd1;
frames[6][21][36] = 8'hb1;
frames[6][21][37] = 8'hb1;
frames[6][21][38] = 8'hb1;
frames[6][21][39] = 8'hb1;
frames[6][22][0] = 8'hac;
frames[6][22][1] = 8'hac;
frames[6][22][2] = 8'hb1;
frames[6][22][3] = 8'hd1;
frames[6][22][4] = 8'hd5;
frames[6][22][5] = 8'hd5;
frames[6][22][6] = 8'hd5;
frames[6][22][7] = 8'hd6;
frames[6][22][8] = 8'hb1;
frames[6][22][9] = 8'hb1;
frames[6][22][10] = 8'h91;
frames[6][22][11] = 8'h91;
frames[6][22][12] = 8'h8d;
frames[6][22][13] = 8'h6d;
frames[6][22][14] = 8'h8d;
frames[6][22][15] = 8'h8d;
frames[6][22][16] = 8'h88;
frames[6][22][17] = 8'h64;
frames[6][22][18] = 8'ha4;
frames[6][22][19] = 8'ha8;
frames[6][22][20] = 8'h8d;
frames[6][22][21] = 8'hb1;
frames[6][22][22] = 8'h91;
frames[6][22][23] = 8'h91;
frames[6][22][24] = 8'h91;
frames[6][22][25] = 8'h91;
frames[6][22][26] = 8'h91;
frames[6][22][27] = 8'hb1;
frames[6][22][28] = 8'h8d;
frames[6][22][29] = 8'h24;
frames[6][22][30] = 8'h8d;
frames[6][22][31] = 8'hb1;
frames[6][22][32] = 8'hb1;
frames[6][22][33] = 8'hb1;
frames[6][22][34] = 8'hb1;
frames[6][22][35] = 8'hb1;
frames[6][22][36] = 8'hb1;
frames[6][22][37] = 8'hb1;
frames[6][22][38] = 8'hb1;
frames[6][22][39] = 8'hb1;
frames[6][23][0] = 8'hac;
frames[6][23][1] = 8'hac;
frames[6][23][2] = 8'hac;
frames[6][23][3] = 8'hb1;
frames[6][23][4] = 8'hb1;
frames[6][23][5] = 8'hd1;
frames[6][23][6] = 8'hd1;
frames[6][23][7] = 8'hd1;
frames[6][23][8] = 8'hb1;
frames[6][23][9] = 8'had;
frames[6][23][10] = 8'h68;
frames[6][23][11] = 8'h8d;
frames[6][23][12] = 8'h8d;
frames[6][23][13] = 8'h8d;
frames[6][23][14] = 8'h8d;
frames[6][23][15] = 8'h8d;
frames[6][23][16] = 8'h89;
frames[6][23][17] = 8'h89;
frames[6][23][18] = 8'h84;
frames[6][23][19] = 8'h84;
frames[6][23][20] = 8'h8d;
frames[6][23][21] = 8'h8d;
frames[6][23][22] = 8'h6d;
frames[6][23][23] = 8'h6d;
frames[6][23][24] = 8'h6d;
frames[6][23][25] = 8'h6d;
frames[6][23][26] = 8'h6d;
frames[6][23][27] = 8'h6d;
frames[6][23][28] = 8'h44;
frames[6][23][29] = 8'h00;
frames[6][23][30] = 8'h8d;
frames[6][23][31] = 8'hb1;
frames[6][23][32] = 8'hd1;
frames[6][23][33] = 8'hb1;
frames[6][23][34] = 8'hb1;
frames[6][23][35] = 8'hb1;
frames[6][23][36] = 8'hb1;
frames[6][23][37] = 8'hb1;
frames[6][23][38] = 8'hb1;
frames[6][23][39] = 8'hb1;
frames[6][24][0] = 8'hac;
frames[6][24][1] = 8'hac;
frames[6][24][2] = 8'hac;
frames[6][24][3] = 8'hac;
frames[6][24][4] = 8'hac;
frames[6][24][5] = 8'hd1;
frames[6][24][6] = 8'hd1;
frames[6][24][7] = 8'hd1;
frames[6][24][8] = 8'hb1;
frames[6][24][9] = 8'hac;
frames[6][24][10] = 8'h20;
frames[6][24][11] = 8'h69;
frames[6][24][12] = 8'h8d;
frames[6][24][13] = 8'h44;
frames[6][24][14] = 8'h44;
frames[6][24][15] = 8'h68;
frames[6][24][16] = 8'h8d;
frames[6][24][17] = 8'h44;
frames[6][24][18] = 8'h44;
frames[6][24][19] = 8'h68;
frames[6][24][20] = 8'h68;
frames[6][24][21] = 8'h69;
frames[6][24][22] = 8'h69;
frames[6][24][23] = 8'h69;
frames[6][24][24] = 8'h69;
frames[6][24][25] = 8'h69;
frames[6][24][26] = 8'h6d;
frames[6][24][27] = 8'h6d;
frames[6][24][28] = 8'h6d;
frames[6][24][29] = 8'h8d;
frames[6][24][30] = 8'hd1;
frames[6][24][31] = 8'hb1;
frames[6][24][32] = 8'hb1;
frames[6][24][33] = 8'hb1;
frames[6][24][34] = 8'hb1;
frames[6][24][35] = 8'hb1;
frames[6][24][36] = 8'hb1;
frames[6][24][37] = 8'hb1;
frames[6][24][38] = 8'hb1;
frames[6][24][39] = 8'hb1;
frames[6][25][0] = 8'h8c;
frames[6][25][1] = 8'hac;
frames[6][25][2] = 8'hac;
frames[6][25][3] = 8'hac;
frames[6][25][4] = 8'hb0;
frames[6][25][5] = 8'hb1;
frames[6][25][6] = 8'hd1;
frames[6][25][7] = 8'hd1;
frames[6][25][8] = 8'hd1;
frames[6][25][9] = 8'hd1;
frames[6][25][10] = 8'h8d;
frames[6][25][11] = 8'hb1;
frames[6][25][12] = 8'h8d;
frames[6][25][13] = 8'h8d;
frames[6][25][14] = 8'h8d;
frames[6][25][15] = 8'h8d;
frames[6][25][16] = 8'hb6;
frames[6][25][17] = 8'h91;
frames[6][25][18] = 8'hb1;
frames[6][25][19] = 8'hb1;
frames[6][25][20] = 8'hb1;
frames[6][25][21] = 8'hb1;
frames[6][25][22] = 8'hd5;
frames[6][25][23] = 8'hd5;
frames[6][25][24] = 8'hd5;
frames[6][25][25] = 8'hd1;
frames[6][25][26] = 8'hd1;
frames[6][25][27] = 8'hd1;
frames[6][25][28] = 8'hd1;
frames[6][25][29] = 8'hb1;
frames[6][25][30] = 8'hb1;
frames[6][25][31] = 8'hb1;
frames[6][25][32] = 8'hb1;
frames[6][25][33] = 8'hb1;
frames[6][25][34] = 8'hb1;
frames[6][25][35] = 8'hb1;
frames[6][25][36] = 8'hb1;
frames[6][25][37] = 8'hb1;
frames[6][25][38] = 8'hb1;
frames[6][25][39] = 8'hb1;
frames[6][26][0] = 8'h8c;
frames[6][26][1] = 8'hac;
frames[6][26][2] = 8'hac;
frames[6][26][3] = 8'hac;
frames[6][26][4] = 8'hac;
frames[6][26][5] = 8'hb1;
frames[6][26][6] = 8'hd1;
frames[6][26][7] = 8'hd1;
frames[6][26][8] = 8'hd1;
frames[6][26][9] = 8'hd1;
frames[6][26][10] = 8'hb1;
frames[6][26][11] = 8'hac;
frames[6][26][12] = 8'had;
frames[6][26][13] = 8'hb1;
frames[6][26][14] = 8'hb1;
frames[6][26][15] = 8'hb1;
frames[6][26][16] = 8'hb1;
frames[6][26][17] = 8'hb1;
frames[6][26][18] = 8'hb1;
frames[6][26][19] = 8'hd6;
frames[6][26][20] = 8'hd6;
frames[6][26][21] = 8'hd6;
frames[6][26][22] = 8'hd6;
frames[6][26][23] = 8'hd6;
frames[6][26][24] = 8'hd1;
frames[6][26][25] = 8'hd1;
frames[6][26][26] = 8'hd1;
frames[6][26][27] = 8'hb1;
frames[6][26][28] = 8'hb1;
frames[6][26][29] = 8'hb1;
frames[6][26][30] = 8'hb1;
frames[6][26][31] = 8'hb1;
frames[6][26][32] = 8'hb1;
frames[6][26][33] = 8'hb1;
frames[6][26][34] = 8'hb1;
frames[6][26][35] = 8'hb1;
frames[6][26][36] = 8'hb1;
frames[6][26][37] = 8'hb1;
frames[6][26][38] = 8'hb1;
frames[6][26][39] = 8'hb1;
frames[6][27][0] = 8'h8c;
frames[6][27][1] = 8'h8c;
frames[6][27][2] = 8'h8c;
frames[6][27][3] = 8'hac;
frames[6][27][4] = 8'hac;
frames[6][27][5] = 8'hb1;
frames[6][27][6] = 8'hb1;
frames[6][27][7] = 8'hb1;
frames[6][27][8] = 8'hd1;
frames[6][27][9] = 8'hd1;
frames[6][27][10] = 8'hb1;
frames[6][27][11] = 8'hb1;
frames[6][27][12] = 8'hb1;
frames[6][27][13] = 8'hb1;
frames[6][27][14] = 8'hb1;
frames[6][27][15] = 8'hb1;
frames[6][27][16] = 8'hac;
frames[6][27][17] = 8'hac;
frames[6][27][18] = 8'hb1;
frames[6][27][19] = 8'hd5;
frames[6][27][20] = 8'hd6;
frames[6][27][21] = 8'hd6;
frames[6][27][22] = 8'hda;
frames[6][27][23] = 8'hd6;
frames[6][27][24] = 8'hd1;
frames[6][27][25] = 8'hb1;
frames[6][27][26] = 8'hb1;
frames[6][27][27] = 8'hb1;
frames[6][27][28] = 8'hb1;
frames[6][27][29] = 8'hb1;
frames[6][27][30] = 8'hb1;
frames[6][27][31] = 8'hb1;
frames[6][27][32] = 8'hb1;
frames[6][27][33] = 8'hb1;
frames[6][27][34] = 8'hb1;
frames[6][27][35] = 8'hb1;
frames[6][27][36] = 8'hb1;
frames[6][27][37] = 8'hb1;
frames[6][27][38] = 8'hb1;
frames[6][27][39] = 8'hb1;
frames[6][28][0] = 8'h88;
frames[6][28][1] = 8'h8c;
frames[6][28][2] = 8'h8c;
frames[6][28][3] = 8'h8c;
frames[6][28][4] = 8'hac;
frames[6][28][5] = 8'hac;
frames[6][28][6] = 8'hb1;
frames[6][28][7] = 8'hb1;
frames[6][28][8] = 8'hd1;
frames[6][28][9] = 8'hd1;
frames[6][28][10] = 8'hb1;
frames[6][28][11] = 8'hb1;
frames[6][28][12] = 8'hb1;
frames[6][28][13] = 8'hb1;
frames[6][28][14] = 8'hb1;
frames[6][28][15] = 8'hb1;
frames[6][28][16] = 8'hac;
frames[6][28][17] = 8'h8c;
frames[6][28][18] = 8'hac;
frames[6][28][19] = 8'had;
frames[6][28][20] = 8'had;
frames[6][28][21] = 8'hb1;
frames[6][28][22] = 8'hd1;
frames[6][28][23] = 8'hd1;
frames[6][28][24] = 8'hb1;
frames[6][28][25] = 8'hb1;
frames[6][28][26] = 8'hb1;
frames[6][28][27] = 8'hb1;
frames[6][28][28] = 8'hb1;
frames[6][28][29] = 8'hb1;
frames[6][28][30] = 8'hb1;
frames[6][28][31] = 8'hb1;
frames[6][28][32] = 8'hb1;
frames[6][28][33] = 8'hb1;
frames[6][28][34] = 8'hb1;
frames[6][28][35] = 8'hb1;
frames[6][28][36] = 8'hb1;
frames[6][28][37] = 8'hb1;
frames[6][28][38] = 8'hb1;
frames[6][28][39] = 8'hb1;
frames[6][29][0] = 8'h88;
frames[6][29][1] = 8'h8c;
frames[6][29][2] = 8'h8c;
frames[6][29][3] = 8'h8c;
frames[6][29][4] = 8'hac;
frames[6][29][5] = 8'hac;
frames[6][29][6] = 8'hac;
frames[6][29][7] = 8'hb1;
frames[6][29][8] = 8'hd1;
frames[6][29][9] = 8'hd1;
frames[6][29][10] = 8'hb1;
frames[6][29][11] = 8'hb1;
frames[6][29][12] = 8'had;
frames[6][29][13] = 8'hb1;
frames[6][29][14] = 8'hb1;
frames[6][29][15] = 8'hb1;
frames[6][29][16] = 8'hac;
frames[6][29][17] = 8'h8c;
frames[6][29][18] = 8'h8c;
frames[6][29][19] = 8'h8c;
frames[6][29][20] = 8'h88;
frames[6][29][21] = 8'h8c;
frames[6][29][22] = 8'had;
frames[6][29][23] = 8'hb1;
frames[6][29][24] = 8'hb1;
frames[6][29][25] = 8'hb1;
frames[6][29][26] = 8'hb1;
frames[6][29][27] = 8'hb1;
frames[6][29][28] = 8'hb1;
frames[6][29][29] = 8'hb1;
frames[6][29][30] = 8'hb1;
frames[6][29][31] = 8'hb1;
frames[6][29][32] = 8'hb1;
frames[6][29][33] = 8'hb1;
frames[6][29][34] = 8'hb1;
frames[6][29][35] = 8'hb1;
frames[6][29][36] = 8'hb1;
frames[6][29][37] = 8'hb1;
frames[6][29][38] = 8'hb1;
frames[6][29][39] = 8'hb1;
frames[7][0][0] = 8'hb1;
frames[7][0][1] = 8'hb1;
frames[7][0][2] = 8'hb1;
frames[7][0][3] = 8'hd1;
frames[7][0][4] = 8'hd1;
frames[7][0][5] = 8'hd1;
frames[7][0][6] = 8'hd1;
frames[7][0][7] = 8'hd5;
frames[7][0][8] = 8'hd1;
frames[7][0][9] = 8'hd1;
frames[7][0][10] = 8'hd1;
frames[7][0][11] = 8'hd5;
frames[7][0][12] = 8'hd5;
frames[7][0][13] = 8'hd5;
frames[7][0][14] = 8'hd5;
frames[7][0][15] = 8'hd5;
frames[7][0][16] = 8'hd5;
frames[7][0][17] = 8'hd1;
frames[7][0][18] = 8'hd5;
frames[7][0][19] = 8'hd1;
frames[7][0][20] = 8'hd1;
frames[7][0][21] = 8'hd1;
frames[7][0][22] = 8'hd5;
frames[7][0][23] = 8'hd5;
frames[7][0][24] = 8'hd5;
frames[7][0][25] = 8'hd5;
frames[7][0][26] = 8'hd5;
frames[7][0][27] = 8'hd1;
frames[7][0][28] = 8'hd1;
frames[7][0][29] = 8'hd1;
frames[7][0][30] = 8'hd1;
frames[7][0][31] = 8'hd1;
frames[7][0][32] = 8'hd1;
frames[7][0][33] = 8'hd5;
frames[7][0][34] = 8'hd1;
frames[7][0][35] = 8'hd1;
frames[7][0][36] = 8'hd1;
frames[7][0][37] = 8'hd1;
frames[7][0][38] = 8'hb1;
frames[7][0][39] = 8'had;
frames[7][1][0] = 8'hb1;
frames[7][1][1] = 8'hb1;
frames[7][1][2] = 8'hb1;
frames[7][1][3] = 8'hd1;
frames[7][1][4] = 8'hd1;
frames[7][1][5] = 8'hd1;
frames[7][1][6] = 8'hd1;
frames[7][1][7] = 8'hd1;
frames[7][1][8] = 8'hd1;
frames[7][1][9] = 8'hd1;
frames[7][1][10] = 8'hd1;
frames[7][1][11] = 8'hd5;
frames[7][1][12] = 8'hd5;
frames[7][1][13] = 8'hd5;
frames[7][1][14] = 8'hd5;
frames[7][1][15] = 8'hd5;
frames[7][1][16] = 8'hd5;
frames[7][1][17] = 8'hd1;
frames[7][1][18] = 8'hd1;
frames[7][1][19] = 8'hd1;
frames[7][1][20] = 8'hd1;
frames[7][1][21] = 8'hd1;
frames[7][1][22] = 8'hd5;
frames[7][1][23] = 8'hd5;
frames[7][1][24] = 8'hd5;
frames[7][1][25] = 8'hd5;
frames[7][1][26] = 8'hd5;
frames[7][1][27] = 8'hd1;
frames[7][1][28] = 8'hd1;
frames[7][1][29] = 8'hd1;
frames[7][1][30] = 8'hd1;
frames[7][1][31] = 8'hd1;
frames[7][1][32] = 8'hd1;
frames[7][1][33] = 8'hd5;
frames[7][1][34] = 8'hd1;
frames[7][1][35] = 8'hd1;
frames[7][1][36] = 8'hd1;
frames[7][1][37] = 8'hd1;
frames[7][1][38] = 8'hb1;
frames[7][1][39] = 8'had;
frames[7][2][0] = 8'hb1;
frames[7][2][1] = 8'hb1;
frames[7][2][2] = 8'hd1;
frames[7][2][3] = 8'hd1;
frames[7][2][4] = 8'hd1;
frames[7][2][5] = 8'hd1;
frames[7][2][6] = 8'hd5;
frames[7][2][7] = 8'hd5;
frames[7][2][8] = 8'hd5;
frames[7][2][9] = 8'hd5;
frames[7][2][10] = 8'hd5;
frames[7][2][11] = 8'hd5;
frames[7][2][12] = 8'hf5;
frames[7][2][13] = 8'hd5;
frames[7][2][14] = 8'hd5;
frames[7][2][15] = 8'hd5;
frames[7][2][16] = 8'hd1;
frames[7][2][17] = 8'hd1;
frames[7][2][18] = 8'hd1;
frames[7][2][19] = 8'hd1;
frames[7][2][20] = 8'hd1;
frames[7][2][21] = 8'hd1;
frames[7][2][22] = 8'hd5;
frames[7][2][23] = 8'hd5;
frames[7][2][24] = 8'hd5;
frames[7][2][25] = 8'hd5;
frames[7][2][26] = 8'hd5;
frames[7][2][27] = 8'hd1;
frames[7][2][28] = 8'hd1;
frames[7][2][29] = 8'hd1;
frames[7][2][30] = 8'hd1;
frames[7][2][31] = 8'hd1;
frames[7][2][32] = 8'hd1;
frames[7][2][33] = 8'hd1;
frames[7][2][34] = 8'hd1;
frames[7][2][35] = 8'hd1;
frames[7][2][36] = 8'hd1;
frames[7][2][37] = 8'hd1;
frames[7][2][38] = 8'hb1;
frames[7][2][39] = 8'hac;
frames[7][3][0] = 8'hb1;
frames[7][3][1] = 8'hb1;
frames[7][3][2] = 8'hd1;
frames[7][3][3] = 8'hd1;
frames[7][3][4] = 8'hd1;
frames[7][3][5] = 8'hd1;
frames[7][3][6] = 8'hd6;
frames[7][3][7] = 8'hd6;
frames[7][3][8] = 8'hd6;
frames[7][3][9] = 8'hd6;
frames[7][3][10] = 8'hd6;
frames[7][3][11] = 8'hd6;
frames[7][3][12] = 8'hf6;
frames[7][3][13] = 8'hd5;
frames[7][3][14] = 8'hd5;
frames[7][3][15] = 8'hd5;
frames[7][3][16] = 8'hd1;
frames[7][3][17] = 8'hd1;
frames[7][3][18] = 8'hd1;
frames[7][3][19] = 8'hd1;
frames[7][3][20] = 8'hd1;
frames[7][3][21] = 8'hd1;
frames[7][3][22] = 8'hd5;
frames[7][3][23] = 8'hd5;
frames[7][3][24] = 8'hd5;
frames[7][3][25] = 8'hd5;
frames[7][3][26] = 8'hd5;
frames[7][3][27] = 8'hd1;
frames[7][3][28] = 8'hd1;
frames[7][3][29] = 8'hd1;
frames[7][3][30] = 8'hd1;
frames[7][3][31] = 8'hd1;
frames[7][3][32] = 8'hd1;
frames[7][3][33] = 8'hd5;
frames[7][3][34] = 8'hd1;
frames[7][3][35] = 8'hd1;
frames[7][3][36] = 8'hd1;
frames[7][3][37] = 8'hd1;
frames[7][3][38] = 8'hb1;
frames[7][3][39] = 8'had;
frames[7][4][0] = 8'hb1;
frames[7][4][1] = 8'hb1;
frames[7][4][2] = 8'hb1;
frames[7][4][3] = 8'hd1;
frames[7][4][4] = 8'hd1;
frames[7][4][5] = 8'hd1;
frames[7][4][6] = 8'hd1;
frames[7][4][7] = 8'hd5;
frames[7][4][8] = 8'hd5;
frames[7][4][9] = 8'hd1;
frames[7][4][10] = 8'hd5;
frames[7][4][11] = 8'hd5;
frames[7][4][12] = 8'hd5;
frames[7][4][13] = 8'hd5;
frames[7][4][14] = 8'hd5;
frames[7][4][15] = 8'hd5;
frames[7][4][16] = 8'hd1;
frames[7][4][17] = 8'hd1;
frames[7][4][18] = 8'hd1;
frames[7][4][19] = 8'hd1;
frames[7][4][20] = 8'hd1;
frames[7][4][21] = 8'hd1;
frames[7][4][22] = 8'hd5;
frames[7][4][23] = 8'hd1;
frames[7][4][24] = 8'hd1;
frames[7][4][25] = 8'hd1;
frames[7][4][26] = 8'hd1;
frames[7][4][27] = 8'hd1;
frames[7][4][28] = 8'hd1;
frames[7][4][29] = 8'hd1;
frames[7][4][30] = 8'hd1;
frames[7][4][31] = 8'hd1;
frames[7][4][32] = 8'hd1;
frames[7][4][33] = 8'hd5;
frames[7][4][34] = 8'hd1;
frames[7][4][35] = 8'hd1;
frames[7][4][36] = 8'hd1;
frames[7][4][37] = 8'hd1;
frames[7][4][38] = 8'hd1;
frames[7][4][39] = 8'had;
frames[7][5][0] = 8'hb1;
frames[7][5][1] = 8'hb1;
frames[7][5][2] = 8'hb1;
frames[7][5][3] = 8'hd1;
frames[7][5][4] = 8'hd1;
frames[7][5][5] = 8'hd1;
frames[7][5][6] = 8'hd1;
frames[7][5][7] = 8'hd1;
frames[7][5][8] = 8'hd1;
frames[7][5][9] = 8'hb1;
frames[7][5][10] = 8'hb1;
frames[7][5][11] = 8'hd1;
frames[7][5][12] = 8'hd5;
frames[7][5][13] = 8'hd5;
frames[7][5][14] = 8'hd1;
frames[7][5][15] = 8'hd5;
frames[7][5][16] = 8'hd1;
frames[7][5][17] = 8'hd1;
frames[7][5][18] = 8'hd1;
frames[7][5][19] = 8'hd1;
frames[7][5][20] = 8'hd1;
frames[7][5][21] = 8'hd1;
frames[7][5][22] = 8'hd1;
frames[7][5][23] = 8'hd1;
frames[7][5][24] = 8'hd1;
frames[7][5][25] = 8'hd1;
frames[7][5][26] = 8'hd1;
frames[7][5][27] = 8'hd1;
frames[7][5][28] = 8'hd1;
frames[7][5][29] = 8'hd1;
frames[7][5][30] = 8'hd5;
frames[7][5][31] = 8'hd5;
frames[7][5][32] = 8'hd5;
frames[7][5][33] = 8'hd5;
frames[7][5][34] = 8'hd5;
frames[7][5][35] = 8'hd5;
frames[7][5][36] = 8'hd1;
frames[7][5][37] = 8'hd1;
frames[7][5][38] = 8'hd1;
frames[7][5][39] = 8'hac;
frames[7][6][0] = 8'hb1;
frames[7][6][1] = 8'hb1;
frames[7][6][2] = 8'hd1;
frames[7][6][3] = 8'hd1;
frames[7][6][4] = 8'hd1;
frames[7][6][5] = 8'hd1;
frames[7][6][6] = 8'hd1;
frames[7][6][7] = 8'hd5;
frames[7][6][8] = 8'hd1;
frames[7][6][9] = 8'hb1;
frames[7][6][10] = 8'hd1;
frames[7][6][11] = 8'hfa;
frames[7][6][12] = 8'hda;
frames[7][6][13] = 8'hda;
frames[7][6][14] = 8'hfa;
frames[7][6][15] = 8'hd5;
frames[7][6][16] = 8'hb1;
frames[7][6][17] = 8'hd6;
frames[7][6][18] = 8'hb1;
frames[7][6][19] = 8'h91;
frames[7][6][20] = 8'h8d;
frames[7][6][21] = 8'hb6;
frames[7][6][22] = 8'hb6;
frames[7][6][23] = 8'h96;
frames[7][6][24] = 8'hb6;
frames[7][6][25] = 8'h96;
frames[7][6][26] = 8'h91;
frames[7][6][27] = 8'h6d;
frames[7][6][28] = 8'h68;
frames[7][6][29] = 8'hd1;
frames[7][6][30] = 8'hd5;
frames[7][6][31] = 8'hd6;
frames[7][6][32] = 8'hd6;
frames[7][6][33] = 8'hd6;
frames[7][6][34] = 8'hd6;
frames[7][6][35] = 8'hd5;
frames[7][6][36] = 8'hd1;
frames[7][6][37] = 8'hd1;
frames[7][6][38] = 8'hd1;
frames[7][6][39] = 8'hac;
frames[7][7][0] = 8'hb1;
frames[7][7][1] = 8'hb1;
frames[7][7][2] = 8'hd1;
frames[7][7][3] = 8'hd1;
frames[7][7][4] = 8'hd1;
frames[7][7][5] = 8'hd1;
frames[7][7][6] = 8'hd1;
frames[7][7][7] = 8'hd1;
frames[7][7][8] = 8'hd1;
frames[7][7][9] = 8'hd1;
frames[7][7][10] = 8'hd6;
frames[7][7][11] = 8'hfe;
frames[7][7][12] = 8'hfe;
frames[7][7][13] = 8'hfe;
frames[7][7][14] = 8'hfe;
frames[7][7][15] = 8'hd6;
frames[7][7][16] = 8'hb1;
frames[7][7][17] = 8'hb1;
frames[7][7][18] = 8'h6d;
frames[7][7][19] = 8'h49;
frames[7][7][20] = 8'h96;
frames[7][7][21] = 8'h96;
frames[7][7][22] = 8'hb6;
frames[7][7][23] = 8'hda;
frames[7][7][24] = 8'hda;
frames[7][7][25] = 8'hb6;
frames[7][7][26] = 8'h92;
frames[7][7][27] = 8'h29;
frames[7][7][28] = 8'h20;
frames[7][7][29] = 8'hb1;
frames[7][7][30] = 8'hd5;
frames[7][7][31] = 8'hd5;
frames[7][7][32] = 8'hd5;
frames[7][7][33] = 8'hd5;
frames[7][7][34] = 8'hd5;
frames[7][7][35] = 8'hd5;
frames[7][7][36] = 8'hd1;
frames[7][7][37] = 8'hd1;
frames[7][7][38] = 8'hd1;
frames[7][7][39] = 8'hac;
frames[7][8][0] = 8'hac;
frames[7][8][1] = 8'hb1;
frames[7][8][2] = 8'hb1;
frames[7][8][3] = 8'hd1;
frames[7][8][4] = 8'hb1;
frames[7][8][5] = 8'hb1;
frames[7][8][6] = 8'hd1;
frames[7][8][7] = 8'hd1;
frames[7][8][8] = 8'hd1;
frames[7][8][9] = 8'hd5;
frames[7][8][10] = 8'hfa;
frames[7][8][11] = 8'hfa;
frames[7][8][12] = 8'hfa;
frames[7][8][13] = 8'hfa;
frames[7][8][14] = 8'hfa;
frames[7][8][15] = 8'hfa;
frames[7][8][16] = 8'hb1;
frames[7][8][17] = 8'h91;
frames[7][8][18] = 8'h6d;
frames[7][8][19] = 8'hb6;
frames[7][8][20] = 8'hb6;
frames[7][8][21] = 8'hda;
frames[7][8][22] = 8'hfa;
frames[7][8][23] = 8'hfa;
frames[7][8][24] = 8'hfa;
frames[7][8][25] = 8'hfa;
frames[7][8][26] = 8'hba;
frames[7][8][27] = 8'h92;
frames[7][8][28] = 8'h44;
frames[7][8][29] = 8'hb1;
frames[7][8][30] = 8'hd1;
frames[7][8][31] = 8'hd5;
frames[7][8][32] = 8'hd1;
frames[7][8][33] = 8'hd5;
frames[7][8][34] = 8'hd5;
frames[7][8][35] = 8'hd5;
frames[7][8][36] = 8'hd1;
frames[7][8][37] = 8'hd1;
frames[7][8][38] = 8'hd1;
frames[7][8][39] = 8'hac;
frames[7][9][0] = 8'hac;
frames[7][9][1] = 8'hb1;
frames[7][9][2] = 8'hb1;
frames[7][9][3] = 8'hd1;
frames[7][9][4] = 8'hb1;
frames[7][9][5] = 8'hb0;
frames[7][9][6] = 8'hd1;
frames[7][9][7] = 8'hd1;
frames[7][9][8] = 8'hb1;
frames[7][9][9] = 8'hb1;
frames[7][9][10] = 8'hd6;
frames[7][9][11] = 8'hfa;
frames[7][9][12] = 8'hfa;
frames[7][9][13] = 8'hfa;
frames[7][9][14] = 8'hfa;
frames[7][9][15] = 8'hfa;
frames[7][9][16] = 8'hb6;
frames[7][9][17] = 8'h91;
frames[7][9][18] = 8'h92;
frames[7][9][19] = 8'hda;
frames[7][9][20] = 8'hfa;
frames[7][9][21] = 8'hfa;
frames[7][9][22] = 8'hfa;
frames[7][9][23] = 8'hfa;
frames[7][9][24] = 8'hfa;
frames[7][9][25] = 8'hfa;
frames[7][9][26] = 8'hfb;
frames[7][9][27] = 8'hda;
frames[7][9][28] = 8'h91;
frames[7][9][29] = 8'hb2;
frames[7][9][30] = 8'hf5;
frames[7][9][31] = 8'hd1;
frames[7][9][32] = 8'hd1;
frames[7][9][33] = 8'hd1;
frames[7][9][34] = 8'hd5;
frames[7][9][35] = 8'hd5;
frames[7][9][36] = 8'hd1;
frames[7][9][37] = 8'hd1;
frames[7][9][38] = 8'hd1;
frames[7][9][39] = 8'hb1;
frames[7][10][0] = 8'hac;
frames[7][10][1] = 8'hb1;
frames[7][10][2] = 8'hb1;
frames[7][10][3] = 8'hb1;
frames[7][10][4] = 8'hb1;
frames[7][10][5] = 8'hb1;
frames[7][10][6] = 8'hd1;
frames[7][10][7] = 8'hd1;
frames[7][10][8] = 8'hb1;
frames[7][10][9] = 8'had;
frames[7][10][10] = 8'hd6;
frames[7][10][11] = 8'hfa;
frames[7][10][12] = 8'hfa;
frames[7][10][13] = 8'hfa;
frames[7][10][14] = 8'hfa;
frames[7][10][15] = 8'hfa;
frames[7][10][16] = 8'hb6;
frames[7][10][17] = 8'h91;
frames[7][10][18] = 8'hd6;
frames[7][10][19] = 8'hff;
frames[7][10][20] = 8'hfa;
frames[7][10][21] = 8'hfa;
frames[7][10][22] = 8'hfa;
frames[7][10][23] = 8'hfa;
frames[7][10][24] = 8'hfa;
frames[7][10][25] = 8'hfa;
frames[7][10][26] = 8'hfb;
frames[7][10][27] = 8'hfb;
frames[7][10][28] = 8'hda;
frames[7][10][29] = 8'hb6;
frames[7][10][30] = 8'hd1;
frames[7][10][31] = 8'hd1;
frames[7][10][32] = 8'hd1;
frames[7][10][33] = 8'hd1;
frames[7][10][34] = 8'hd5;
frames[7][10][35] = 8'hd5;
frames[7][10][36] = 8'hd1;
frames[7][10][37] = 8'hb1;
frames[7][10][38] = 8'hb1;
frames[7][10][39] = 8'hb1;
frames[7][11][0] = 8'hac;
frames[7][11][1] = 8'hb0;
frames[7][11][2] = 8'hb1;
frames[7][11][3] = 8'hb1;
frames[7][11][4] = 8'hb1;
frames[7][11][5] = 8'hb1;
frames[7][11][6] = 8'hd1;
frames[7][11][7] = 8'hd1;
frames[7][11][8] = 8'hb1;
frames[7][11][9] = 8'had;
frames[7][11][10] = 8'hd5;
frames[7][11][11] = 8'hda;
frames[7][11][12] = 8'hda;
frames[7][11][13] = 8'hfa;
frames[7][11][14] = 8'hfa;
frames[7][11][15] = 8'hfa;
frames[7][11][16] = 8'hb2;
frames[7][11][17] = 8'hb2;
frames[7][11][18] = 8'hfa;
frames[7][11][19] = 8'hff;
frames[7][11][20] = 8'hfa;
frames[7][11][21] = 8'hfa;
frames[7][11][22] = 8'hfa;
frames[7][11][23] = 8'hfa;
frames[7][11][24] = 8'hfa;
frames[7][11][25] = 8'hfa;
frames[7][11][26] = 8'hfa;
frames[7][11][27] = 8'hfa;
frames[7][11][28] = 8'hda;
frames[7][11][29] = 8'hb6;
frames[7][11][30] = 8'hd1;
frames[7][11][31] = 8'hd1;
frames[7][11][32] = 8'hd1;
frames[7][11][33] = 8'hd1;
frames[7][11][34] = 8'hd5;
frames[7][11][35] = 8'hd5;
frames[7][11][36] = 8'hd1;
frames[7][11][37] = 8'hb1;
frames[7][11][38] = 8'hb1;
frames[7][11][39] = 8'hb1;
frames[7][12][0] = 8'hac;
frames[7][12][1] = 8'had;
frames[7][12][2] = 8'hb1;
frames[7][12][3] = 8'hb1;
frames[7][12][4] = 8'hb1;
frames[7][12][5] = 8'hb1;
frames[7][12][6] = 8'hd1;
frames[7][12][7] = 8'hd1;
frames[7][12][8] = 8'hb1;
frames[7][12][9] = 8'hac;
frames[7][12][10] = 8'hb1;
frames[7][12][11] = 8'hd6;
frames[7][12][12] = 8'hfa;
frames[7][12][13] = 8'hfa;
frames[7][12][14] = 8'hfa;
frames[7][12][15] = 8'hd6;
frames[7][12][16] = 8'hb1;
frames[7][12][17] = 8'hb6;
frames[7][12][18] = 8'hfb;
frames[7][12][19] = 8'hfb;
frames[7][12][20] = 8'hfb;
frames[7][12][21] = 8'hfa;
frames[7][12][22] = 8'hfa;
frames[7][12][23] = 8'hfa;
frames[7][12][24] = 8'hfa;
frames[7][12][25] = 8'hfa;
frames[7][12][26] = 8'hfa;
frames[7][12][27] = 8'hfa;
frames[7][12][28] = 8'hfa;
frames[7][12][29] = 8'hb6;
frames[7][12][30] = 8'hd1;
frames[7][12][31] = 8'hd1;
frames[7][12][32] = 8'hd1;
frames[7][12][33] = 8'hd1;
frames[7][12][34] = 8'hd5;
frames[7][12][35] = 8'hd5;
frames[7][12][36] = 8'hd1;
frames[7][12][37] = 8'hb1;
frames[7][12][38] = 8'hb1;
frames[7][12][39] = 8'hb1;
frames[7][13][0] = 8'hac;
frames[7][13][1] = 8'hac;
frames[7][13][2] = 8'hb1;
frames[7][13][3] = 8'hb0;
frames[7][13][4] = 8'hb0;
frames[7][13][5] = 8'hb1;
frames[7][13][6] = 8'hb1;
frames[7][13][7] = 8'hb1;
frames[7][13][8] = 8'had;
frames[7][13][9] = 8'hac;
frames[7][13][10] = 8'h8d;
frames[7][13][11] = 8'hb1;
frames[7][13][12] = 8'hd6;
frames[7][13][13] = 8'hfa;
frames[7][13][14] = 8'hda;
frames[7][13][15] = 8'hb1;
frames[7][13][16] = 8'h91;
frames[7][13][17] = 8'hb6;
frames[7][13][18] = 8'hfa;
frames[7][13][19] = 8'hff;
frames[7][13][20] = 8'hfb;
frames[7][13][21] = 8'hfb;
frames[7][13][22] = 8'hfa;
frames[7][13][23] = 8'hfa;
frames[7][13][24] = 8'hfa;
frames[7][13][25] = 8'hfa;
frames[7][13][26] = 8'hfa;
frames[7][13][27] = 8'hfa;
frames[7][13][28] = 8'hfa;
frames[7][13][29] = 8'hb6;
frames[7][13][30] = 8'hd1;
frames[7][13][31] = 8'hd1;
frames[7][13][32] = 8'hd1;
frames[7][13][33] = 8'hd1;
frames[7][13][34] = 8'hd5;
frames[7][13][35] = 8'hd5;
frames[7][13][36] = 8'hd1;
frames[7][13][37] = 8'hb1;
frames[7][13][38] = 8'hb1;
frames[7][13][39] = 8'hb1;
frames[7][14][0] = 8'hac;
frames[7][14][1] = 8'hac;
frames[7][14][2] = 8'hb1;
frames[7][14][3] = 8'hb1;
frames[7][14][4] = 8'hb0;
frames[7][14][5] = 8'hb1;
frames[7][14][6] = 8'hb1;
frames[7][14][7] = 8'hac;
frames[7][14][8] = 8'hac;
frames[7][14][9] = 8'hac;
frames[7][14][10] = 8'h8d;
frames[7][14][11] = 8'h91;
frames[7][14][12] = 8'hb1;
frames[7][14][13] = 8'hb5;
frames[7][14][14] = 8'h91;
frames[7][14][15] = 8'hb1;
frames[7][14][16] = 8'h91;
frames[7][14][17] = 8'h91;
frames[7][14][18] = 8'hfa;
frames[7][14][19] = 8'hff;
frames[7][14][20] = 8'hfb;
frames[7][14][21] = 8'hfa;
frames[7][14][22] = 8'hfa;
frames[7][14][23] = 8'hfa;
frames[7][14][24] = 8'hfa;
frames[7][14][25] = 8'hfa;
frames[7][14][26] = 8'hfa;
frames[7][14][27] = 8'hfa;
frames[7][14][28] = 8'hfa;
frames[7][14][29] = 8'hb6;
frames[7][14][30] = 8'hd1;
frames[7][14][31] = 8'hd1;
frames[7][14][32] = 8'hd1;
frames[7][14][33] = 8'hd1;
frames[7][14][34] = 8'hd1;
frames[7][14][35] = 8'hd5;
frames[7][14][36] = 8'hd1;
frames[7][14][37] = 8'hb1;
frames[7][14][38] = 8'hb1;
frames[7][14][39] = 8'hb1;
frames[7][15][0] = 8'hac;
frames[7][15][1] = 8'hac;
frames[7][15][2] = 8'hac;
frames[7][15][3] = 8'hac;
frames[7][15][4] = 8'hac;
frames[7][15][5] = 8'hb1;
frames[7][15][6] = 8'hb1;
frames[7][15][7] = 8'hac;
frames[7][15][8] = 8'hac;
frames[7][15][9] = 8'hac;
frames[7][15][10] = 8'h89;
frames[7][15][11] = 8'h89;
frames[7][15][12] = 8'h89;
frames[7][15][13] = 8'h8d;
frames[7][15][14] = 8'h91;
frames[7][15][15] = 8'hb1;
frames[7][15][16] = 8'h8d;
frames[7][15][17] = 8'h8d;
frames[7][15][18] = 8'hfa;
frames[7][15][19] = 8'hff;
frames[7][15][20] = 8'hff;
frames[7][15][21] = 8'hfb;
frames[7][15][22] = 8'hfa;
frames[7][15][23] = 8'hfa;
frames[7][15][24] = 8'hfa;
frames[7][15][25] = 8'hfa;
frames[7][15][26] = 8'hfa;
frames[7][15][27] = 8'hfa;
frames[7][15][28] = 8'hda;
frames[7][15][29] = 8'hb6;
frames[7][15][30] = 8'hd1;
frames[7][15][31] = 8'hd1;
frames[7][15][32] = 8'hd1;
frames[7][15][33] = 8'hd1;
frames[7][15][34] = 8'hd1;
frames[7][15][35] = 8'hd5;
frames[7][15][36] = 8'hd1;
frames[7][15][37] = 8'hb1;
frames[7][15][38] = 8'hb1;
frames[7][15][39] = 8'hb1;
frames[7][16][0] = 8'hac;
frames[7][16][1] = 8'hac;
frames[7][16][2] = 8'hac;
frames[7][16][3] = 8'hac;
frames[7][16][4] = 8'hac;
frames[7][16][5] = 8'hb0;
frames[7][16][6] = 8'hb1;
frames[7][16][7] = 8'hac;
frames[7][16][8] = 8'hac;
frames[7][16][9] = 8'hac;
frames[7][16][10] = 8'had;
frames[7][16][11] = 8'h64;
frames[7][16][12] = 8'h60;
frames[7][16][13] = 8'h84;
frames[7][16][14] = 8'h8d;
frames[7][16][15] = 8'hb1;
frames[7][16][16] = 8'h91;
frames[7][16][17] = 8'h8d;
frames[7][16][18] = 8'hd6;
frames[7][16][19] = 8'hff;
frames[7][16][20] = 8'hfa;
frames[7][16][21] = 8'hfa;
frames[7][16][22] = 8'hfa;
frames[7][16][23] = 8'hfa;
frames[7][16][24] = 8'hfa;
frames[7][16][25] = 8'hfa;
frames[7][16][26] = 8'hfa;
frames[7][16][27] = 8'hfa;
frames[7][16][28] = 8'hda;
frames[7][16][29] = 8'h91;
frames[7][16][30] = 8'hb1;
frames[7][16][31] = 8'hd1;
frames[7][16][32] = 8'hd1;
frames[7][16][33] = 8'hd1;
frames[7][16][34] = 8'hd1;
frames[7][16][35] = 8'hd5;
frames[7][16][36] = 8'hd1;
frames[7][16][37] = 8'hb1;
frames[7][16][38] = 8'hb1;
frames[7][16][39] = 8'hb1;
frames[7][17][0] = 8'hac;
frames[7][17][1] = 8'hac;
frames[7][17][2] = 8'hac;
frames[7][17][3] = 8'hac;
frames[7][17][4] = 8'hb0;
frames[7][17][5] = 8'hb1;
frames[7][17][6] = 8'hb0;
frames[7][17][7] = 8'hac;
frames[7][17][8] = 8'hac;
frames[7][17][9] = 8'h8c;
frames[7][17][10] = 8'h84;
frames[7][17][11] = 8'h60;
frames[7][17][12] = 8'h60;
frames[7][17][13] = 8'h60;
frames[7][17][14] = 8'h69;
frames[7][17][15] = 8'h8d;
frames[7][17][16] = 8'h91;
frames[7][17][17] = 8'h8d;
frames[7][17][18] = 8'hb1;
frames[7][17][19] = 8'hfb;
frames[7][17][20] = 8'hfb;
frames[7][17][21] = 8'hfa;
frames[7][17][22] = 8'hfa;
frames[7][17][23] = 8'hfa;
frames[7][17][24] = 8'hfa;
frames[7][17][25] = 8'hfa;
frames[7][17][26] = 8'hfa;
frames[7][17][27] = 8'hfa;
frames[7][17][28] = 8'hb6;
frames[7][17][29] = 8'h6d;
frames[7][17][30] = 8'hb1;
frames[7][17][31] = 8'hd1;
frames[7][17][32] = 8'hd1;
frames[7][17][33] = 8'hd1;
frames[7][17][34] = 8'hd1;
frames[7][17][35] = 8'hd1;
frames[7][17][36] = 8'hd1;
frames[7][17][37] = 8'hb1;
frames[7][17][38] = 8'hb1;
frames[7][17][39] = 8'hb1;
frames[7][18][0] = 8'hac;
frames[7][18][1] = 8'hac;
frames[7][18][2] = 8'hac;
frames[7][18][3] = 8'hac;
frames[7][18][4] = 8'hb0;
frames[7][18][5] = 8'hd1;
frames[7][18][6] = 8'hd1;
frames[7][18][7] = 8'hb1;
frames[7][18][8] = 8'hac;
frames[7][18][9] = 8'h8c;
frames[7][18][10] = 8'h64;
frames[7][18][11] = 8'h60;
frames[7][18][12] = 8'h60;
frames[7][18][13] = 8'h60;
frames[7][18][14] = 8'h68;
frames[7][18][15] = 8'h8d;
frames[7][18][16] = 8'h8d;
frames[7][18][17] = 8'h8d;
frames[7][18][18] = 8'h6d;
frames[7][18][19] = 8'hd6;
frames[7][18][20] = 8'hfa;
frames[7][18][21] = 8'hfb;
frames[7][18][22] = 8'hfa;
frames[7][18][23] = 8'hfa;
frames[7][18][24] = 8'hfa;
frames[7][18][25] = 8'hfa;
frames[7][18][26] = 8'hfa;
frames[7][18][27] = 8'hda;
frames[7][18][28] = 8'hb6;
frames[7][18][29] = 8'h48;
frames[7][18][30] = 8'hb1;
frames[7][18][31] = 8'hb1;
frames[7][18][32] = 8'hd1;
frames[7][18][33] = 8'hd1;
frames[7][18][34] = 8'hd1;
frames[7][18][35] = 8'hd1;
frames[7][18][36] = 8'hd1;
frames[7][18][37] = 8'hb1;
frames[7][18][38] = 8'hb1;
frames[7][18][39] = 8'hb1;
frames[7][19][0] = 8'hac;
frames[7][19][1] = 8'hac;
frames[7][19][2] = 8'hac;
frames[7][19][3] = 8'hac;
frames[7][19][4] = 8'hb0;
frames[7][19][5] = 8'hd1;
frames[7][19][6] = 8'hd1;
frames[7][19][7] = 8'hd1;
frames[7][19][8] = 8'hac;
frames[7][19][9] = 8'h8c;
frames[7][19][10] = 8'h84;
frames[7][19][11] = 8'h40;
frames[7][19][12] = 8'h60;
frames[7][19][13] = 8'h60;
frames[7][19][14] = 8'h69;
frames[7][19][15] = 8'h8d;
frames[7][19][16] = 8'h8d;
frames[7][19][17] = 8'h69;
frames[7][19][18] = 8'h68;
frames[7][19][19] = 8'h8d;
frames[7][19][20] = 8'hda;
frames[7][19][21] = 8'hdb;
frames[7][19][22] = 8'hfa;
frames[7][19][23] = 8'hda;
frames[7][19][24] = 8'hda;
frames[7][19][25] = 8'hda;
frames[7][19][26] = 8'hda;
frames[7][19][27] = 8'hb6;
frames[7][19][28] = 8'h8d;
frames[7][19][29] = 8'h44;
frames[7][19][30] = 8'hb1;
frames[7][19][31] = 8'hb1;
frames[7][19][32] = 8'hd1;
frames[7][19][33] = 8'hd1;
frames[7][19][34] = 8'hd1;
frames[7][19][35] = 8'hd1;
frames[7][19][36] = 8'hd1;
frames[7][19][37] = 8'hb1;
frames[7][19][38] = 8'hb1;
frames[7][19][39] = 8'hb1;
frames[7][20][0] = 8'hac;
frames[7][20][1] = 8'hac;
frames[7][20][2] = 8'hac;
frames[7][20][3] = 8'hac;
frames[7][20][4] = 8'hac;
frames[7][20][5] = 8'hb1;
frames[7][20][6] = 8'hd1;
frames[7][20][7] = 8'hb1;
frames[7][20][8] = 8'hac;
frames[7][20][9] = 8'had;
frames[7][20][10] = 8'h89;
frames[7][20][11] = 8'h64;
frames[7][20][12] = 8'h64;
frames[7][20][13] = 8'h88;
frames[7][20][14] = 8'h69;
frames[7][20][15] = 8'h8d;
frames[7][20][16] = 8'ha9;
frames[7][20][17] = 8'h88;
frames[7][20][18] = 8'ha8;
frames[7][20][19] = 8'ha4;
frames[7][20][20] = 8'h92;
frames[7][20][21] = 8'hba;
frames[7][20][22] = 8'hb6;
frames[7][20][23] = 8'h96;
frames[7][20][24] = 8'hb6;
frames[7][20][25] = 8'hba;
frames[7][20][26] = 8'hb6;
frames[7][20][27] = 8'hb6;
frames[7][20][28] = 8'h8d;
frames[7][20][29] = 8'h44;
frames[7][20][30] = 8'hb1;
frames[7][20][31] = 8'hb1;
frames[7][20][32] = 8'hd1;
frames[7][20][33] = 8'hd1;
frames[7][20][34] = 8'hb1;
frames[7][20][35] = 8'hd1;
frames[7][20][36] = 8'hb1;
frames[7][20][37] = 8'hb1;
frames[7][20][38] = 8'hb1;
frames[7][20][39] = 8'hb1;
frames[7][21][0] = 8'hac;
frames[7][21][1] = 8'hac;
frames[7][21][2] = 8'hb1;
frames[7][21][3] = 8'hd1;
frames[7][21][4] = 8'hd1;
frames[7][21][5] = 8'hd1;
frames[7][21][6] = 8'hd5;
frames[7][21][7] = 8'hd5;
frames[7][21][8] = 8'hb1;
frames[7][21][9] = 8'hb1;
frames[7][21][10] = 8'h8d;
frames[7][21][11] = 8'h8d;
frames[7][21][12] = 8'h91;
frames[7][21][13] = 8'h8d;
frames[7][21][14] = 8'h8d;
frames[7][21][15] = 8'h8d;
frames[7][21][16] = 8'ha8;
frames[7][21][17] = 8'h64;
frames[7][21][18] = 8'ha8;
frames[7][21][19] = 8'ha4;
frames[7][21][20] = 8'h8d;
frames[7][21][21] = 8'hb1;
frames[7][21][22] = 8'hb6;
frames[7][21][23] = 8'hb6;
frames[7][21][24] = 8'hb6;
frames[7][21][25] = 8'hb6;
frames[7][21][26] = 8'hb2;
frames[7][21][27] = 8'hb2;
frames[7][21][28] = 8'h91;
frames[7][21][29] = 8'h44;
frames[7][21][30] = 8'had;
frames[7][21][31] = 8'hb1;
frames[7][21][32] = 8'hd1;
frames[7][21][33] = 8'hd1;
frames[7][21][34] = 8'hb1;
frames[7][21][35] = 8'hd1;
frames[7][21][36] = 8'hb1;
frames[7][21][37] = 8'hb1;
frames[7][21][38] = 8'hb1;
frames[7][21][39] = 8'hb1;
frames[7][22][0] = 8'hac;
frames[7][22][1] = 8'hac;
frames[7][22][2] = 8'hb1;
frames[7][22][3] = 8'hd5;
frames[7][22][4] = 8'hd5;
frames[7][22][5] = 8'hd5;
frames[7][22][6] = 8'hd5;
frames[7][22][7] = 8'hd6;
frames[7][22][8] = 8'hb1;
frames[7][22][9] = 8'hb1;
frames[7][22][10] = 8'h91;
frames[7][22][11] = 8'h91;
frames[7][22][12] = 8'h8d;
frames[7][22][13] = 8'h6d;
frames[7][22][14] = 8'h8d;
frames[7][22][15] = 8'h8d;
frames[7][22][16] = 8'h88;
frames[7][22][17] = 8'h64;
frames[7][22][18] = 8'ha4;
frames[7][22][19] = 8'ha8;
frames[7][22][20] = 8'h8d;
frames[7][22][21] = 8'hb1;
frames[7][22][22] = 8'h91;
frames[7][22][23] = 8'h91;
frames[7][22][24] = 8'h91;
frames[7][22][25] = 8'h91;
frames[7][22][26] = 8'h91;
frames[7][22][27] = 8'hb1;
frames[7][22][28] = 8'h91;
frames[7][22][29] = 8'h24;
frames[7][22][30] = 8'h8c;
frames[7][22][31] = 8'hb1;
frames[7][22][32] = 8'hb1;
frames[7][22][33] = 8'hb1;
frames[7][22][34] = 8'hb1;
frames[7][22][35] = 8'hb1;
frames[7][22][36] = 8'hb1;
frames[7][22][37] = 8'hb1;
frames[7][22][38] = 8'hb1;
frames[7][22][39] = 8'hb1;
frames[7][23][0] = 8'hac;
frames[7][23][1] = 8'hac;
frames[7][23][2] = 8'hac;
frames[7][23][3] = 8'hb1;
frames[7][23][4] = 8'hb1;
frames[7][23][5] = 8'hd1;
frames[7][23][6] = 8'hd1;
frames[7][23][7] = 8'hd1;
frames[7][23][8] = 8'hb1;
frames[7][23][9] = 8'had;
frames[7][23][10] = 8'h68;
frames[7][23][11] = 8'h8d;
frames[7][23][12] = 8'h8d;
frames[7][23][13] = 8'h8d;
frames[7][23][14] = 8'h8d;
frames[7][23][15] = 8'h8d;
frames[7][23][16] = 8'h89;
frames[7][23][17] = 8'h89;
frames[7][23][18] = 8'h84;
frames[7][23][19] = 8'h84;
frames[7][23][20] = 8'h8d;
frames[7][23][21] = 8'h8d;
frames[7][23][22] = 8'h6d;
frames[7][23][23] = 8'h6d;
frames[7][23][24] = 8'h6d;
frames[7][23][25] = 8'h6d;
frames[7][23][26] = 8'h6d;
frames[7][23][27] = 8'h6d;
frames[7][23][28] = 8'h44;
frames[7][23][29] = 8'h00;
frames[7][23][30] = 8'h8d;
frames[7][23][31] = 8'hb1;
frames[7][23][32] = 8'hb1;
frames[7][23][33] = 8'hb1;
frames[7][23][34] = 8'hb1;
frames[7][23][35] = 8'hb1;
frames[7][23][36] = 8'hb1;
frames[7][23][37] = 8'hb1;
frames[7][23][38] = 8'hb1;
frames[7][23][39] = 8'hb1;
frames[7][24][0] = 8'hac;
frames[7][24][1] = 8'hac;
frames[7][24][2] = 8'hac;
frames[7][24][3] = 8'hac;
frames[7][24][4] = 8'hac;
frames[7][24][5] = 8'hd1;
frames[7][24][6] = 8'hd1;
frames[7][24][7] = 8'hd1;
frames[7][24][8] = 8'hb1;
frames[7][24][9] = 8'hac;
frames[7][24][10] = 8'h20;
frames[7][24][11] = 8'h69;
frames[7][24][12] = 8'h8d;
frames[7][24][13] = 8'h44;
frames[7][24][14] = 8'h44;
frames[7][24][15] = 8'h68;
frames[7][24][16] = 8'h8d;
frames[7][24][17] = 8'h44;
frames[7][24][18] = 8'h44;
frames[7][24][19] = 8'h68;
frames[7][24][20] = 8'h68;
frames[7][24][21] = 8'h69;
frames[7][24][22] = 8'h69;
frames[7][24][23] = 8'h69;
frames[7][24][24] = 8'h69;
frames[7][24][25] = 8'h69;
frames[7][24][26] = 8'h6d;
frames[7][24][27] = 8'h6d;
frames[7][24][28] = 8'h6d;
frames[7][24][29] = 8'h8d;
frames[7][24][30] = 8'hb1;
frames[7][24][31] = 8'hb1;
frames[7][24][32] = 8'hb1;
frames[7][24][33] = 8'hb1;
frames[7][24][34] = 8'hb1;
frames[7][24][35] = 8'hb1;
frames[7][24][36] = 8'hb1;
frames[7][24][37] = 8'hb1;
frames[7][24][38] = 8'hb1;
frames[7][24][39] = 8'hb1;
frames[7][25][0] = 8'hac;
frames[7][25][1] = 8'hac;
frames[7][25][2] = 8'hac;
frames[7][25][3] = 8'hac;
frames[7][25][4] = 8'hb0;
frames[7][25][5] = 8'hb1;
frames[7][25][6] = 8'hd1;
frames[7][25][7] = 8'hd1;
frames[7][25][8] = 8'hd1;
frames[7][25][9] = 8'hd1;
frames[7][25][10] = 8'h8d;
frames[7][25][11] = 8'hb1;
frames[7][25][12] = 8'h8d;
frames[7][25][13] = 8'h8d;
frames[7][25][14] = 8'h8d;
frames[7][25][15] = 8'h8d;
frames[7][25][16] = 8'hb6;
frames[7][25][17] = 8'hb1;
frames[7][25][18] = 8'hb1;
frames[7][25][19] = 8'hb1;
frames[7][25][20] = 8'hb1;
frames[7][25][21] = 8'hb1;
frames[7][25][22] = 8'hd5;
frames[7][25][23] = 8'hd5;
frames[7][25][24] = 8'hd1;
frames[7][25][25] = 8'hd1;
frames[7][25][26] = 8'hd1;
frames[7][25][27] = 8'hd1;
frames[7][25][28] = 8'hd1;
frames[7][25][29] = 8'hd1;
frames[7][25][30] = 8'hb1;
frames[7][25][31] = 8'hb1;
frames[7][25][32] = 8'hb1;
frames[7][25][33] = 8'hb1;
frames[7][25][34] = 8'hb1;
frames[7][25][35] = 8'hb1;
frames[7][25][36] = 8'hb1;
frames[7][25][37] = 8'hb1;
frames[7][25][38] = 8'hb1;
frames[7][25][39] = 8'hb1;
frames[7][26][0] = 8'h8c;
frames[7][26][1] = 8'hac;
frames[7][26][2] = 8'hac;
frames[7][26][3] = 8'hac;
frames[7][26][4] = 8'hac;
frames[7][26][5] = 8'hb1;
frames[7][26][6] = 8'hd1;
frames[7][26][7] = 8'hd1;
frames[7][26][8] = 8'hd1;
frames[7][26][9] = 8'hd1;
frames[7][26][10] = 8'hd1;
frames[7][26][11] = 8'hac;
frames[7][26][12] = 8'had;
frames[7][26][13] = 8'hb1;
frames[7][26][14] = 8'hb1;
frames[7][26][15] = 8'hb1;
frames[7][26][16] = 8'hb1;
frames[7][26][17] = 8'hb1;
frames[7][26][18] = 8'hb1;
frames[7][26][19] = 8'hd6;
frames[7][26][20] = 8'hd6;
frames[7][26][21] = 8'hd6;
frames[7][26][22] = 8'hd6;
frames[7][26][23] = 8'hd6;
frames[7][26][24] = 8'hd1;
frames[7][26][25] = 8'hd1;
frames[7][26][26] = 8'hd1;
frames[7][26][27] = 8'hb1;
frames[7][26][28] = 8'hb1;
frames[7][26][29] = 8'hb1;
frames[7][26][30] = 8'hb1;
frames[7][26][31] = 8'hb1;
frames[7][26][32] = 8'hb1;
frames[7][26][33] = 8'hb1;
frames[7][26][34] = 8'hb1;
frames[7][26][35] = 8'hb1;
frames[7][26][36] = 8'hb1;
frames[7][26][37] = 8'hb1;
frames[7][26][38] = 8'hb1;
frames[7][26][39] = 8'hb1;
frames[7][27][0] = 8'h8c;
frames[7][27][1] = 8'h8c;
frames[7][27][2] = 8'hac;
frames[7][27][3] = 8'hac;
frames[7][27][4] = 8'hac;
frames[7][27][5] = 8'hb1;
frames[7][27][6] = 8'hd1;
frames[7][27][7] = 8'hd1;
frames[7][27][8] = 8'hd1;
frames[7][27][9] = 8'hd1;
frames[7][27][10] = 8'hb1;
frames[7][27][11] = 8'hb1;
frames[7][27][12] = 8'hb1;
frames[7][27][13] = 8'hb1;
frames[7][27][14] = 8'hb1;
frames[7][27][15] = 8'hb1;
frames[7][27][16] = 8'hac;
frames[7][27][17] = 8'hac;
frames[7][27][18] = 8'hb1;
frames[7][27][19] = 8'hd5;
frames[7][27][20] = 8'hd6;
frames[7][27][21] = 8'hd6;
frames[7][27][22] = 8'hda;
frames[7][27][23] = 8'hd6;
frames[7][27][24] = 8'hd1;
frames[7][27][25] = 8'hb1;
frames[7][27][26] = 8'hb1;
frames[7][27][27] = 8'hb1;
frames[7][27][28] = 8'hb1;
frames[7][27][29] = 8'hb1;
frames[7][27][30] = 8'hb1;
frames[7][27][31] = 8'hb1;
frames[7][27][32] = 8'hb1;
frames[7][27][33] = 8'hb1;
frames[7][27][34] = 8'hb1;
frames[7][27][35] = 8'hb1;
frames[7][27][36] = 8'hb1;
frames[7][27][37] = 8'hb1;
frames[7][27][38] = 8'hb1;
frames[7][27][39] = 8'hb1;
frames[7][28][0] = 8'h88;
frames[7][28][1] = 8'h8c;
frames[7][28][2] = 8'h8c;
frames[7][28][3] = 8'h8c;
frames[7][28][4] = 8'hac;
frames[7][28][5] = 8'hac;
frames[7][28][6] = 8'hb1;
frames[7][28][7] = 8'hb1;
frames[7][28][8] = 8'hd1;
frames[7][28][9] = 8'hd1;
frames[7][28][10] = 8'hb1;
frames[7][28][11] = 8'hb1;
frames[7][28][12] = 8'hb1;
frames[7][28][13] = 8'hb1;
frames[7][28][14] = 8'hb1;
frames[7][28][15] = 8'hb1;
frames[7][28][16] = 8'hac;
frames[7][28][17] = 8'h8c;
frames[7][28][18] = 8'hac;
frames[7][28][19] = 8'had;
frames[7][28][20] = 8'had;
frames[7][28][21] = 8'hb1;
frames[7][28][22] = 8'hd5;
frames[7][28][23] = 8'hd5;
frames[7][28][24] = 8'hb1;
frames[7][28][25] = 8'hb1;
frames[7][28][26] = 8'hb1;
frames[7][28][27] = 8'hb1;
frames[7][28][28] = 8'hb1;
frames[7][28][29] = 8'hb1;
frames[7][28][30] = 8'hb1;
frames[7][28][31] = 8'hb1;
frames[7][28][32] = 8'hb1;
frames[7][28][33] = 8'hb1;
frames[7][28][34] = 8'hb1;
frames[7][28][35] = 8'hb1;
frames[7][28][36] = 8'hb1;
frames[7][28][37] = 8'hb1;
frames[7][28][38] = 8'hb1;
frames[7][28][39] = 8'had;
frames[7][29][0] = 8'h88;
frames[7][29][1] = 8'h8c;
frames[7][29][2] = 8'h8c;
frames[7][29][3] = 8'h8c;
frames[7][29][4] = 8'hac;
frames[7][29][5] = 8'hac;
frames[7][29][6] = 8'hac;
frames[7][29][7] = 8'hb1;
frames[7][29][8] = 8'hd1;
frames[7][29][9] = 8'hb1;
frames[7][29][10] = 8'hb1;
frames[7][29][11] = 8'hb1;
frames[7][29][12] = 8'had;
frames[7][29][13] = 8'hb1;
frames[7][29][14] = 8'hb1;
frames[7][29][15] = 8'hb1;
frames[7][29][16] = 8'hac;
frames[7][29][17] = 8'h8c;
frames[7][29][18] = 8'h8c;
frames[7][29][19] = 8'h8c;
frames[7][29][20] = 8'h88;
frames[7][29][21] = 8'h8c;
frames[7][29][22] = 8'had;
frames[7][29][23] = 8'hb1;
frames[7][29][24] = 8'hb1;
frames[7][29][25] = 8'hb1;
frames[7][29][26] = 8'hb1;
frames[7][29][27] = 8'hb1;
frames[7][29][28] = 8'hb1;
frames[7][29][29] = 8'hb1;
frames[7][29][30] = 8'hb1;
frames[7][29][31] = 8'hb1;
frames[7][29][32] = 8'hb1;
frames[7][29][33] = 8'hb1;
frames[7][29][34] = 8'hb1;
frames[7][29][35] = 8'hb1;
frames[7][29][36] = 8'hb1;
frames[7][29][37] = 8'hb1;
frames[7][29][38] = 8'hb1;
frames[7][29][39] = 8'hb1;
frames[8][0][0] = 8'hb1;
frames[8][0][1] = 8'hb1;
frames[8][0][2] = 8'hb1;
frames[8][0][3] = 8'hd1;
frames[8][0][4] = 8'hd1;
frames[8][0][5] = 8'hd1;
frames[8][0][6] = 8'hd1;
frames[8][0][7] = 8'hd5;
frames[8][0][8] = 8'hd1;
frames[8][0][9] = 8'hd1;
frames[8][0][10] = 8'hd1;
frames[8][0][11] = 8'hd5;
frames[8][0][12] = 8'hd5;
frames[8][0][13] = 8'hd5;
frames[8][0][14] = 8'hd5;
frames[8][0][15] = 8'hd5;
frames[8][0][16] = 8'hd5;
frames[8][0][17] = 8'hd1;
frames[8][0][18] = 8'hd5;
frames[8][0][19] = 8'hd1;
frames[8][0][20] = 8'hd1;
frames[8][0][21] = 8'hd1;
frames[8][0][22] = 8'hd5;
frames[8][0][23] = 8'hd5;
frames[8][0][24] = 8'hd5;
frames[8][0][25] = 8'hd5;
frames[8][0][26] = 8'hd5;
frames[8][0][27] = 8'hd1;
frames[8][0][28] = 8'hd1;
frames[8][0][29] = 8'hd1;
frames[8][0][30] = 8'hd1;
frames[8][0][31] = 8'hd1;
frames[8][0][32] = 8'hd1;
frames[8][0][33] = 8'hd5;
frames[8][0][34] = 8'hd1;
frames[8][0][35] = 8'hd1;
frames[8][0][36] = 8'hd1;
frames[8][0][37] = 8'hd1;
frames[8][0][38] = 8'hb1;
frames[8][0][39] = 8'had;
frames[8][1][0] = 8'hb1;
frames[8][1][1] = 8'hb1;
frames[8][1][2] = 8'hb1;
frames[8][1][3] = 8'hd1;
frames[8][1][4] = 8'hd1;
frames[8][1][5] = 8'hd1;
frames[8][1][6] = 8'hd1;
frames[8][1][7] = 8'hd1;
frames[8][1][8] = 8'hd1;
frames[8][1][9] = 8'hd1;
frames[8][1][10] = 8'hd1;
frames[8][1][11] = 8'hd5;
frames[8][1][12] = 8'hd5;
frames[8][1][13] = 8'hd5;
frames[8][1][14] = 8'hd5;
frames[8][1][15] = 8'hd5;
frames[8][1][16] = 8'hd5;
frames[8][1][17] = 8'hd1;
frames[8][1][18] = 8'hd1;
frames[8][1][19] = 8'hd1;
frames[8][1][20] = 8'hd1;
frames[8][1][21] = 8'hd1;
frames[8][1][22] = 8'hd5;
frames[8][1][23] = 8'hd5;
frames[8][1][24] = 8'hd5;
frames[8][1][25] = 8'hd5;
frames[8][1][26] = 8'hd5;
frames[8][1][27] = 8'hd1;
frames[8][1][28] = 8'hd1;
frames[8][1][29] = 8'hd1;
frames[8][1][30] = 8'hd1;
frames[8][1][31] = 8'hd1;
frames[8][1][32] = 8'hd1;
frames[8][1][33] = 8'hd5;
frames[8][1][34] = 8'hd1;
frames[8][1][35] = 8'hd1;
frames[8][1][36] = 8'hd1;
frames[8][1][37] = 8'hd1;
frames[8][1][38] = 8'hb1;
frames[8][1][39] = 8'had;
frames[8][2][0] = 8'hb1;
frames[8][2][1] = 8'hb1;
frames[8][2][2] = 8'hd1;
frames[8][2][3] = 8'hd1;
frames[8][2][4] = 8'hd1;
frames[8][2][5] = 8'hd1;
frames[8][2][6] = 8'hd5;
frames[8][2][7] = 8'hd5;
frames[8][2][8] = 8'hd5;
frames[8][2][9] = 8'hd5;
frames[8][2][10] = 8'hd5;
frames[8][2][11] = 8'hd5;
frames[8][2][12] = 8'hf5;
frames[8][2][13] = 8'hd5;
frames[8][2][14] = 8'hd5;
frames[8][2][15] = 8'hd5;
frames[8][2][16] = 8'hd1;
frames[8][2][17] = 8'hd1;
frames[8][2][18] = 8'hd1;
frames[8][2][19] = 8'hd1;
frames[8][2][20] = 8'hd1;
frames[8][2][21] = 8'hd1;
frames[8][2][22] = 8'hd5;
frames[8][2][23] = 8'hd5;
frames[8][2][24] = 8'hd5;
frames[8][2][25] = 8'hd5;
frames[8][2][26] = 8'hd5;
frames[8][2][27] = 8'hd1;
frames[8][2][28] = 8'hd1;
frames[8][2][29] = 8'hd1;
frames[8][2][30] = 8'hd1;
frames[8][2][31] = 8'hd1;
frames[8][2][32] = 8'hd1;
frames[8][2][33] = 8'hd5;
frames[8][2][34] = 8'hd1;
frames[8][2][35] = 8'hd1;
frames[8][2][36] = 8'hd1;
frames[8][2][37] = 8'hd1;
frames[8][2][38] = 8'hb1;
frames[8][2][39] = 8'hac;
frames[8][3][0] = 8'hb1;
frames[8][3][1] = 8'hb1;
frames[8][3][2] = 8'hd1;
frames[8][3][3] = 8'hd1;
frames[8][3][4] = 8'hd1;
frames[8][3][5] = 8'hd1;
frames[8][3][6] = 8'hd6;
frames[8][3][7] = 8'hd6;
frames[8][3][8] = 8'hd6;
frames[8][3][9] = 8'hd6;
frames[8][3][10] = 8'hd6;
frames[8][3][11] = 8'hd6;
frames[8][3][12] = 8'hf6;
frames[8][3][13] = 8'hd5;
frames[8][3][14] = 8'hd5;
frames[8][3][15] = 8'hd5;
frames[8][3][16] = 8'hd1;
frames[8][3][17] = 8'hd1;
frames[8][3][18] = 8'hd1;
frames[8][3][19] = 8'hd1;
frames[8][3][20] = 8'hd1;
frames[8][3][21] = 8'hd1;
frames[8][3][22] = 8'hd5;
frames[8][3][23] = 8'hd5;
frames[8][3][24] = 8'hd5;
frames[8][3][25] = 8'hd5;
frames[8][3][26] = 8'hd5;
frames[8][3][27] = 8'hd1;
frames[8][3][28] = 8'hd1;
frames[8][3][29] = 8'hd1;
frames[8][3][30] = 8'hd1;
frames[8][3][31] = 8'hd1;
frames[8][3][32] = 8'hd1;
frames[8][3][33] = 8'hd5;
frames[8][3][34] = 8'hd1;
frames[8][3][35] = 8'hd1;
frames[8][3][36] = 8'hd1;
frames[8][3][37] = 8'hd1;
frames[8][3][38] = 8'hb1;
frames[8][3][39] = 8'had;
frames[8][4][0] = 8'hb1;
frames[8][4][1] = 8'hb1;
frames[8][4][2] = 8'hd1;
frames[8][4][3] = 8'hd1;
frames[8][4][4] = 8'hd1;
frames[8][4][5] = 8'hd1;
frames[8][4][6] = 8'hd1;
frames[8][4][7] = 8'hd5;
frames[8][4][8] = 8'hd5;
frames[8][4][9] = 8'hd1;
frames[8][4][10] = 8'hd5;
frames[8][4][11] = 8'hd5;
frames[8][4][12] = 8'hd5;
frames[8][4][13] = 8'hd5;
frames[8][4][14] = 8'hd5;
frames[8][4][15] = 8'hd5;
frames[8][4][16] = 8'hd1;
frames[8][4][17] = 8'hd1;
frames[8][4][18] = 8'hd1;
frames[8][4][19] = 8'hd1;
frames[8][4][20] = 8'hd1;
frames[8][4][21] = 8'hd1;
frames[8][4][22] = 8'hd5;
frames[8][4][23] = 8'hd1;
frames[8][4][24] = 8'hd1;
frames[8][4][25] = 8'hd1;
frames[8][4][26] = 8'hd1;
frames[8][4][27] = 8'hd1;
frames[8][4][28] = 8'hd1;
frames[8][4][29] = 8'hd1;
frames[8][4][30] = 8'hd1;
frames[8][4][31] = 8'hd1;
frames[8][4][32] = 8'hd1;
frames[8][4][33] = 8'hd5;
frames[8][4][34] = 8'hd1;
frames[8][4][35] = 8'hd1;
frames[8][4][36] = 8'hd1;
frames[8][4][37] = 8'hd1;
frames[8][4][38] = 8'hd1;
frames[8][4][39] = 8'had;
frames[8][5][0] = 8'hb1;
frames[8][5][1] = 8'hb1;
frames[8][5][2] = 8'hb1;
frames[8][5][3] = 8'hd1;
frames[8][5][4] = 8'hd1;
frames[8][5][5] = 8'hd1;
frames[8][5][6] = 8'hd1;
frames[8][5][7] = 8'hd1;
frames[8][5][8] = 8'hd1;
frames[8][5][9] = 8'hb1;
frames[8][5][10] = 8'hd1;
frames[8][5][11] = 8'hd1;
frames[8][5][12] = 8'hd5;
frames[8][5][13] = 8'hd5;
frames[8][5][14] = 8'hd1;
frames[8][5][15] = 8'hd5;
frames[8][5][16] = 8'hd1;
frames[8][5][17] = 8'hd1;
frames[8][5][18] = 8'hd1;
frames[8][5][19] = 8'hd1;
frames[8][5][20] = 8'hd1;
frames[8][5][21] = 8'hd1;
frames[8][5][22] = 8'hd1;
frames[8][5][23] = 8'hd1;
frames[8][5][24] = 8'hd1;
frames[8][5][25] = 8'hd1;
frames[8][5][26] = 8'hd1;
frames[8][5][27] = 8'hd1;
frames[8][5][28] = 8'hd1;
frames[8][5][29] = 8'hd1;
frames[8][5][30] = 8'hd5;
frames[8][5][31] = 8'hd5;
frames[8][5][32] = 8'hd5;
frames[8][5][33] = 8'hd5;
frames[8][5][34] = 8'hd5;
frames[8][5][35] = 8'hd5;
frames[8][5][36] = 8'hd1;
frames[8][5][37] = 8'hd1;
frames[8][5][38] = 8'hd1;
frames[8][5][39] = 8'hac;
frames[8][6][0] = 8'hb1;
frames[8][6][1] = 8'hb1;
frames[8][6][2] = 8'hd1;
frames[8][6][3] = 8'hd1;
frames[8][6][4] = 8'hd1;
frames[8][6][5] = 8'hd1;
frames[8][6][6] = 8'hd1;
frames[8][6][7] = 8'hd5;
frames[8][6][8] = 8'hd1;
frames[8][6][9] = 8'hb1;
frames[8][6][10] = 8'hd1;
frames[8][6][11] = 8'hfa;
frames[8][6][12] = 8'hda;
frames[8][6][13] = 8'hda;
frames[8][6][14] = 8'hfa;
frames[8][6][15] = 8'hd5;
frames[8][6][16] = 8'hb1;
frames[8][6][17] = 8'hd6;
frames[8][6][18] = 8'hb1;
frames[8][6][19] = 8'h91;
frames[8][6][20] = 8'h8d;
frames[8][6][21] = 8'hb6;
frames[8][6][22] = 8'hb6;
frames[8][6][23] = 8'h96;
frames[8][6][24] = 8'hb6;
frames[8][6][25] = 8'h96;
frames[8][6][26] = 8'h91;
frames[8][6][27] = 8'h6d;
frames[8][6][28] = 8'h68;
frames[8][6][29] = 8'hd1;
frames[8][6][30] = 8'hd5;
frames[8][6][31] = 8'hd6;
frames[8][6][32] = 8'hd6;
frames[8][6][33] = 8'hd6;
frames[8][6][34] = 8'hd6;
frames[8][6][35] = 8'hd5;
frames[8][6][36] = 8'hd1;
frames[8][6][37] = 8'hd1;
frames[8][6][38] = 8'hd1;
frames[8][6][39] = 8'hac;
frames[8][7][0] = 8'hb1;
frames[8][7][1] = 8'hb1;
frames[8][7][2] = 8'hd1;
frames[8][7][3] = 8'hd1;
frames[8][7][4] = 8'hd1;
frames[8][7][5] = 8'hb1;
frames[8][7][6] = 8'hd1;
frames[8][7][7] = 8'hd1;
frames[8][7][8] = 8'hd1;
frames[8][7][9] = 8'hb1;
frames[8][7][10] = 8'hd6;
frames[8][7][11] = 8'hfe;
frames[8][7][12] = 8'hfe;
frames[8][7][13] = 8'hfe;
frames[8][7][14] = 8'hfe;
frames[8][7][15] = 8'hd6;
frames[8][7][16] = 8'hb1;
frames[8][7][17] = 8'hb1;
frames[8][7][18] = 8'h8d;
frames[8][7][19] = 8'h49;
frames[8][7][20] = 8'h96;
frames[8][7][21] = 8'h96;
frames[8][7][22] = 8'hb6;
frames[8][7][23] = 8'hda;
frames[8][7][24] = 8'hda;
frames[8][7][25] = 8'hb6;
frames[8][7][26] = 8'h92;
frames[8][7][27] = 8'h29;
frames[8][7][28] = 8'h20;
frames[8][7][29] = 8'hb1;
frames[8][7][30] = 8'hd5;
frames[8][7][31] = 8'hd5;
frames[8][7][32] = 8'hd5;
frames[8][7][33] = 8'hd5;
frames[8][7][34] = 8'hd5;
frames[8][7][35] = 8'hd5;
frames[8][7][36] = 8'hd1;
frames[8][7][37] = 8'hd1;
frames[8][7][38] = 8'hd1;
frames[8][7][39] = 8'hac;
frames[8][8][0] = 8'hac;
frames[8][8][1] = 8'hb1;
frames[8][8][2] = 8'hb1;
frames[8][8][3] = 8'hd1;
frames[8][8][4] = 8'hb1;
frames[8][8][5] = 8'hb1;
frames[8][8][6] = 8'hd1;
frames[8][8][7] = 8'hd1;
frames[8][8][8] = 8'hd1;
frames[8][8][9] = 8'hd5;
frames[8][8][10] = 8'hfa;
frames[8][8][11] = 8'hfa;
frames[8][8][12] = 8'hfa;
frames[8][8][13] = 8'hfa;
frames[8][8][14] = 8'hfa;
frames[8][8][15] = 8'hfa;
frames[8][8][16] = 8'hb1;
frames[8][8][17] = 8'h91;
frames[8][8][18] = 8'h6d;
frames[8][8][19] = 8'hb6;
frames[8][8][20] = 8'hb6;
frames[8][8][21] = 8'hda;
frames[8][8][22] = 8'hfa;
frames[8][8][23] = 8'hfa;
frames[8][8][24] = 8'hfa;
frames[8][8][25] = 8'hfa;
frames[8][8][26] = 8'hba;
frames[8][8][27] = 8'h92;
frames[8][8][28] = 8'h44;
frames[8][8][29] = 8'hb1;
frames[8][8][30] = 8'hd1;
frames[8][8][31] = 8'hd5;
frames[8][8][32] = 8'hd1;
frames[8][8][33] = 8'hd5;
frames[8][8][34] = 8'hd5;
frames[8][8][35] = 8'hd5;
frames[8][8][36] = 8'hd1;
frames[8][8][37] = 8'hd1;
frames[8][8][38] = 8'hd1;
frames[8][8][39] = 8'hac;
frames[8][9][0] = 8'hac;
frames[8][9][1] = 8'hb1;
frames[8][9][2] = 8'hb1;
frames[8][9][3] = 8'hd1;
frames[8][9][4] = 8'hb1;
frames[8][9][5] = 8'hb1;
frames[8][9][6] = 8'hd1;
frames[8][9][7] = 8'hd1;
frames[8][9][8] = 8'hb1;
frames[8][9][9] = 8'hb1;
frames[8][9][10] = 8'hd6;
frames[8][9][11] = 8'hfa;
frames[8][9][12] = 8'hfa;
frames[8][9][13] = 8'hfa;
frames[8][9][14] = 8'hfa;
frames[8][9][15] = 8'hfa;
frames[8][9][16] = 8'hb6;
frames[8][9][17] = 8'h91;
frames[8][9][18] = 8'h92;
frames[8][9][19] = 8'hda;
frames[8][9][20] = 8'hfa;
frames[8][9][21] = 8'hfa;
frames[8][9][22] = 8'hfa;
frames[8][9][23] = 8'hfa;
frames[8][9][24] = 8'hfa;
frames[8][9][25] = 8'hfa;
frames[8][9][26] = 8'hfb;
frames[8][9][27] = 8'hda;
frames[8][9][28] = 8'h91;
frames[8][9][29] = 8'hb2;
frames[8][9][30] = 8'hf5;
frames[8][9][31] = 8'hd1;
frames[8][9][32] = 8'hd1;
frames[8][9][33] = 8'hd1;
frames[8][9][34] = 8'hd5;
frames[8][9][35] = 8'hd5;
frames[8][9][36] = 8'hd1;
frames[8][9][37] = 8'hd1;
frames[8][9][38] = 8'hd1;
frames[8][9][39] = 8'hb1;
frames[8][10][0] = 8'hac;
frames[8][10][1] = 8'hb1;
frames[8][10][2] = 8'hb1;
frames[8][10][3] = 8'hd1;
frames[8][10][4] = 8'hb1;
frames[8][10][5] = 8'hb1;
frames[8][10][6] = 8'hd1;
frames[8][10][7] = 8'hd1;
frames[8][10][8] = 8'hb1;
frames[8][10][9] = 8'had;
frames[8][10][10] = 8'hd6;
frames[8][10][11] = 8'hfa;
frames[8][10][12] = 8'hfa;
frames[8][10][13] = 8'hfa;
frames[8][10][14] = 8'hfa;
frames[8][10][15] = 8'hfa;
frames[8][10][16] = 8'hb6;
frames[8][10][17] = 8'h91;
frames[8][10][18] = 8'hd6;
frames[8][10][19] = 8'hff;
frames[8][10][20] = 8'hfa;
frames[8][10][21] = 8'hfa;
frames[8][10][22] = 8'hfa;
frames[8][10][23] = 8'hfa;
frames[8][10][24] = 8'hfa;
frames[8][10][25] = 8'hfa;
frames[8][10][26] = 8'hfb;
frames[8][10][27] = 8'hfb;
frames[8][10][28] = 8'hda;
frames[8][10][29] = 8'hb6;
frames[8][10][30] = 8'hd1;
frames[8][10][31] = 8'hd1;
frames[8][10][32] = 8'hd1;
frames[8][10][33] = 8'hd1;
frames[8][10][34] = 8'hd5;
frames[8][10][35] = 8'hd5;
frames[8][10][36] = 8'hd1;
frames[8][10][37] = 8'hb1;
frames[8][10][38] = 8'hd1;
frames[8][10][39] = 8'hb1;
frames[8][11][0] = 8'hac;
frames[8][11][1] = 8'hac;
frames[8][11][2] = 8'hb1;
frames[8][11][3] = 8'hb1;
frames[8][11][4] = 8'hb1;
frames[8][11][5] = 8'hb1;
frames[8][11][6] = 8'hd1;
frames[8][11][7] = 8'hd1;
frames[8][11][8] = 8'hb1;
frames[8][11][9] = 8'had;
frames[8][11][10] = 8'hd5;
frames[8][11][11] = 8'hda;
frames[8][11][12] = 8'hda;
frames[8][11][13] = 8'hfa;
frames[8][11][14] = 8'hfa;
frames[8][11][15] = 8'hfa;
frames[8][11][16] = 8'hb2;
frames[8][11][17] = 8'hb2;
frames[8][11][18] = 8'hfa;
frames[8][11][19] = 8'hff;
frames[8][11][20] = 8'hfa;
frames[8][11][21] = 8'hfa;
frames[8][11][22] = 8'hfa;
frames[8][11][23] = 8'hfa;
frames[8][11][24] = 8'hfa;
frames[8][11][25] = 8'hfa;
frames[8][11][26] = 8'hfa;
frames[8][11][27] = 8'hfa;
frames[8][11][28] = 8'hda;
frames[8][11][29] = 8'hb6;
frames[8][11][30] = 8'hd1;
frames[8][11][31] = 8'hd1;
frames[8][11][32] = 8'hd1;
frames[8][11][33] = 8'hd1;
frames[8][11][34] = 8'hd5;
frames[8][11][35] = 8'hd5;
frames[8][11][36] = 8'hd1;
frames[8][11][37] = 8'hb1;
frames[8][11][38] = 8'hb1;
frames[8][11][39] = 8'hb1;
frames[8][12][0] = 8'hac;
frames[8][12][1] = 8'hac;
frames[8][12][2] = 8'hb1;
frames[8][12][3] = 8'hb0;
frames[8][12][4] = 8'hb1;
frames[8][12][5] = 8'hb1;
frames[8][12][6] = 8'hd1;
frames[8][12][7] = 8'hb1;
frames[8][12][8] = 8'hb1;
frames[8][12][9] = 8'hac;
frames[8][12][10] = 8'hb1;
frames[8][12][11] = 8'hd6;
frames[8][12][12] = 8'hfa;
frames[8][12][13] = 8'hfa;
frames[8][12][14] = 8'hfa;
frames[8][12][15] = 8'hd6;
frames[8][12][16] = 8'hb1;
frames[8][12][17] = 8'hb6;
frames[8][12][18] = 8'hfb;
frames[8][12][19] = 8'hfb;
frames[8][12][20] = 8'hfb;
frames[8][12][21] = 8'hfa;
frames[8][12][22] = 8'hfa;
frames[8][12][23] = 8'hfa;
frames[8][12][24] = 8'hfa;
frames[8][12][25] = 8'hfa;
frames[8][12][26] = 8'hfa;
frames[8][12][27] = 8'hfa;
frames[8][12][28] = 8'hfa;
frames[8][12][29] = 8'hb6;
frames[8][12][30] = 8'hd1;
frames[8][12][31] = 8'hd1;
frames[8][12][32] = 8'hd1;
frames[8][12][33] = 8'hd1;
frames[8][12][34] = 8'hd5;
frames[8][12][35] = 8'hd5;
frames[8][12][36] = 8'hd1;
frames[8][12][37] = 8'hb1;
frames[8][12][38] = 8'hb1;
frames[8][12][39] = 8'hb1;
frames[8][13][0] = 8'hac;
frames[8][13][1] = 8'hac;
frames[8][13][2] = 8'hb1;
frames[8][13][3] = 8'hb1;
frames[8][13][4] = 8'hb1;
frames[8][13][5] = 8'hb1;
frames[8][13][6] = 8'hb1;
frames[8][13][7] = 8'hb1;
frames[8][13][8] = 8'had;
frames[8][13][9] = 8'hac;
frames[8][13][10] = 8'h8d;
frames[8][13][11] = 8'hb1;
frames[8][13][12] = 8'hd6;
frames[8][13][13] = 8'hfa;
frames[8][13][14] = 8'hda;
frames[8][13][15] = 8'hb1;
frames[8][13][16] = 8'h91;
frames[8][13][17] = 8'hb6;
frames[8][13][18] = 8'hfa;
frames[8][13][19] = 8'hff;
frames[8][13][20] = 8'hfb;
frames[8][13][21] = 8'hfb;
frames[8][13][22] = 8'hfa;
frames[8][13][23] = 8'hfa;
frames[8][13][24] = 8'hfa;
frames[8][13][25] = 8'hfa;
frames[8][13][26] = 8'hfa;
frames[8][13][27] = 8'hfa;
frames[8][13][28] = 8'hfa;
frames[8][13][29] = 8'hb6;
frames[8][13][30] = 8'hd1;
frames[8][13][31] = 8'hd1;
frames[8][13][32] = 8'hd1;
frames[8][13][33] = 8'hd1;
frames[8][13][34] = 8'hd5;
frames[8][13][35] = 8'hd5;
frames[8][13][36] = 8'hd1;
frames[8][13][37] = 8'hb1;
frames[8][13][38] = 8'hb1;
frames[8][13][39] = 8'hb1;
frames[8][14][0] = 8'hac;
frames[8][14][1] = 8'hac;
frames[8][14][2] = 8'hb1;
frames[8][14][3] = 8'hb1;
frames[8][14][4] = 8'hb1;
frames[8][14][5] = 8'hb1;
frames[8][14][6] = 8'hb1;
frames[8][14][7] = 8'hac;
frames[8][14][8] = 8'hac;
frames[8][14][9] = 8'hac;
frames[8][14][10] = 8'h8d;
frames[8][14][11] = 8'h91;
frames[8][14][12] = 8'hb1;
frames[8][14][13] = 8'hb5;
frames[8][14][14] = 8'h91;
frames[8][14][15] = 8'hb1;
frames[8][14][16] = 8'h91;
frames[8][14][17] = 8'h91;
frames[8][14][18] = 8'hfa;
frames[8][14][19] = 8'hff;
frames[8][14][20] = 8'hfb;
frames[8][14][21] = 8'hfa;
frames[8][14][22] = 8'hfa;
frames[8][14][23] = 8'hfa;
frames[8][14][24] = 8'hfa;
frames[8][14][25] = 8'hfa;
frames[8][14][26] = 8'hfa;
frames[8][14][27] = 8'hfa;
frames[8][14][28] = 8'hfa;
frames[8][14][29] = 8'hb6;
frames[8][14][30] = 8'hd1;
frames[8][14][31] = 8'hd1;
frames[8][14][32] = 8'hd1;
frames[8][14][33] = 8'hd1;
frames[8][14][34] = 8'hd1;
frames[8][14][35] = 8'hd5;
frames[8][14][36] = 8'hd1;
frames[8][14][37] = 8'hb1;
frames[8][14][38] = 8'hb1;
frames[8][14][39] = 8'hb1;
frames[8][15][0] = 8'hac;
frames[8][15][1] = 8'hac;
frames[8][15][2] = 8'hac;
frames[8][15][3] = 8'hac;
frames[8][15][4] = 8'hac;
frames[8][15][5] = 8'hb1;
frames[8][15][6] = 8'hb1;
frames[8][15][7] = 8'hac;
frames[8][15][8] = 8'hac;
frames[8][15][9] = 8'hac;
frames[8][15][10] = 8'h89;
frames[8][15][11] = 8'h89;
frames[8][15][12] = 8'h88;
frames[8][15][13] = 8'h8d;
frames[8][15][14] = 8'h91;
frames[8][15][15] = 8'h91;
frames[8][15][16] = 8'h8d;
frames[8][15][17] = 8'h8d;
frames[8][15][18] = 8'hfa;
frames[8][15][19] = 8'hff;
frames[8][15][20] = 8'hff;
frames[8][15][21] = 8'hfa;
frames[8][15][22] = 8'hfa;
frames[8][15][23] = 8'hfa;
frames[8][15][24] = 8'hfa;
frames[8][15][25] = 8'hfa;
frames[8][15][26] = 8'hfa;
frames[8][15][27] = 8'hfa;
frames[8][15][28] = 8'hda;
frames[8][15][29] = 8'hb6;
frames[8][15][30] = 8'hd1;
frames[8][15][31] = 8'hd1;
frames[8][15][32] = 8'hd1;
frames[8][15][33] = 8'hd1;
frames[8][15][34] = 8'hd1;
frames[8][15][35] = 8'hd5;
frames[8][15][36] = 8'hd1;
frames[8][15][37] = 8'hb1;
frames[8][15][38] = 8'hb1;
frames[8][15][39] = 8'hb1;
frames[8][16][0] = 8'hac;
frames[8][16][1] = 8'hac;
frames[8][16][2] = 8'hac;
frames[8][16][3] = 8'hac;
frames[8][16][4] = 8'hac;
frames[8][16][5] = 8'hb0;
frames[8][16][6] = 8'hb1;
frames[8][16][7] = 8'hac;
frames[8][16][8] = 8'hac;
frames[8][16][9] = 8'hac;
frames[8][16][10] = 8'had;
frames[8][16][11] = 8'h64;
frames[8][16][12] = 8'h60;
frames[8][16][13] = 8'h84;
frames[8][16][14] = 8'h8d;
frames[8][16][15] = 8'hb1;
frames[8][16][16] = 8'h91;
frames[8][16][17] = 8'h8d;
frames[8][16][18] = 8'hd6;
frames[8][16][19] = 8'hff;
frames[8][16][20] = 8'hfa;
frames[8][16][21] = 8'hfa;
frames[8][16][22] = 8'hfa;
frames[8][16][23] = 8'hfa;
frames[8][16][24] = 8'hfa;
frames[8][16][25] = 8'hfa;
frames[8][16][26] = 8'hfa;
frames[8][16][27] = 8'hfa;
frames[8][16][28] = 8'hda;
frames[8][16][29] = 8'h91;
frames[8][16][30] = 8'hb1;
frames[8][16][31] = 8'hd1;
frames[8][16][32] = 8'hd1;
frames[8][16][33] = 8'hd1;
frames[8][16][34] = 8'hd1;
frames[8][16][35] = 8'hd5;
frames[8][16][36] = 8'hd1;
frames[8][16][37] = 8'hb1;
frames[8][16][38] = 8'hb1;
frames[8][16][39] = 8'hb1;
frames[8][17][0] = 8'hac;
frames[8][17][1] = 8'hac;
frames[8][17][2] = 8'hac;
frames[8][17][3] = 8'hac;
frames[8][17][4] = 8'hb0;
frames[8][17][5] = 8'hb1;
frames[8][17][6] = 8'hb1;
frames[8][17][7] = 8'hac;
frames[8][17][8] = 8'hac;
frames[8][17][9] = 8'h8c;
frames[8][17][10] = 8'h84;
frames[8][17][11] = 8'h60;
frames[8][17][12] = 8'h60;
frames[8][17][13] = 8'h60;
frames[8][17][14] = 8'h69;
frames[8][17][15] = 8'h8d;
frames[8][17][16] = 8'h91;
frames[8][17][17] = 8'h8d;
frames[8][17][18] = 8'hb1;
frames[8][17][19] = 8'hfb;
frames[8][17][20] = 8'hfb;
frames[8][17][21] = 8'hfa;
frames[8][17][22] = 8'hfa;
frames[8][17][23] = 8'hfa;
frames[8][17][24] = 8'hfa;
frames[8][17][25] = 8'hfa;
frames[8][17][26] = 8'hfa;
frames[8][17][27] = 8'hfa;
frames[8][17][28] = 8'hb6;
frames[8][17][29] = 8'h6d;
frames[8][17][30] = 8'hb1;
frames[8][17][31] = 8'hd1;
frames[8][17][32] = 8'hd1;
frames[8][17][33] = 8'hd1;
frames[8][17][34] = 8'hd1;
frames[8][17][35] = 8'hd1;
frames[8][17][36] = 8'hd1;
frames[8][17][37] = 8'hb1;
frames[8][17][38] = 8'hb1;
frames[8][17][39] = 8'hb1;
frames[8][18][0] = 8'hac;
frames[8][18][1] = 8'hac;
frames[8][18][2] = 8'hac;
frames[8][18][3] = 8'hac;
frames[8][18][4] = 8'hb0;
frames[8][18][5] = 8'hd1;
frames[8][18][6] = 8'hd1;
frames[8][18][7] = 8'hb1;
frames[8][18][8] = 8'hac;
frames[8][18][9] = 8'h8c;
frames[8][18][10] = 8'h64;
frames[8][18][11] = 8'h60;
frames[8][18][12] = 8'h60;
frames[8][18][13] = 8'h60;
frames[8][18][14] = 8'h68;
frames[8][18][15] = 8'h8d;
frames[8][18][16] = 8'h8d;
frames[8][18][17] = 8'h8d;
frames[8][18][18] = 8'h6d;
frames[8][18][19] = 8'hd6;
frames[8][18][20] = 8'hfa;
frames[8][18][21] = 8'hfb;
frames[8][18][22] = 8'hfa;
frames[8][18][23] = 8'hfa;
frames[8][18][24] = 8'hfa;
frames[8][18][25] = 8'hfa;
frames[8][18][26] = 8'hfa;
frames[8][18][27] = 8'hda;
frames[8][18][28] = 8'hb6;
frames[8][18][29] = 8'h48;
frames[8][18][30] = 8'hb1;
frames[8][18][31] = 8'hb1;
frames[8][18][32] = 8'hd1;
frames[8][18][33] = 8'hd1;
frames[8][18][34] = 8'hd1;
frames[8][18][35] = 8'hd1;
frames[8][18][36] = 8'hd1;
frames[8][18][37] = 8'hb1;
frames[8][18][38] = 8'hb1;
frames[8][18][39] = 8'hb1;
frames[8][19][0] = 8'hac;
frames[8][19][1] = 8'hac;
frames[8][19][2] = 8'hac;
frames[8][19][3] = 8'hac;
frames[8][19][4] = 8'hb0;
frames[8][19][5] = 8'hd1;
frames[8][19][6] = 8'hd1;
frames[8][19][7] = 8'hd1;
frames[8][19][8] = 8'hac;
frames[8][19][9] = 8'h8c;
frames[8][19][10] = 8'h84;
frames[8][19][11] = 8'h40;
frames[8][19][12] = 8'h60;
frames[8][19][13] = 8'h60;
frames[8][19][14] = 8'h69;
frames[8][19][15] = 8'h8d;
frames[8][19][16] = 8'h8d;
frames[8][19][17] = 8'h69;
frames[8][19][18] = 8'h68;
frames[8][19][19] = 8'h8d;
frames[8][19][20] = 8'hda;
frames[8][19][21] = 8'hdb;
frames[8][19][22] = 8'hfa;
frames[8][19][23] = 8'hda;
frames[8][19][24] = 8'hda;
frames[8][19][25] = 8'hda;
frames[8][19][26] = 8'hda;
frames[8][19][27] = 8'hb6;
frames[8][19][28] = 8'h8d;
frames[8][19][29] = 8'h44;
frames[8][19][30] = 8'hb1;
frames[8][19][31] = 8'hb1;
frames[8][19][32] = 8'hd1;
frames[8][19][33] = 8'hd1;
frames[8][19][34] = 8'hd1;
frames[8][19][35] = 8'hd1;
frames[8][19][36] = 8'hd1;
frames[8][19][37] = 8'hb1;
frames[8][19][38] = 8'hb1;
frames[8][19][39] = 8'hb1;
frames[8][20][0] = 8'hac;
frames[8][20][1] = 8'hac;
frames[8][20][2] = 8'hac;
frames[8][20][3] = 8'hac;
frames[8][20][4] = 8'hb0;
frames[8][20][5] = 8'hb1;
frames[8][20][6] = 8'hd1;
frames[8][20][7] = 8'hb1;
frames[8][20][8] = 8'hac;
frames[8][20][9] = 8'had;
frames[8][20][10] = 8'h89;
frames[8][20][11] = 8'h64;
frames[8][20][12] = 8'h64;
frames[8][20][13] = 8'h88;
frames[8][20][14] = 8'h69;
frames[8][20][15] = 8'h8d;
frames[8][20][16] = 8'ha9;
frames[8][20][17] = 8'h84;
frames[8][20][18] = 8'ha8;
frames[8][20][19] = 8'ha4;
frames[8][20][20] = 8'h92;
frames[8][20][21] = 8'hba;
frames[8][20][22] = 8'hb6;
frames[8][20][23] = 8'h96;
frames[8][20][24] = 8'hb6;
frames[8][20][25] = 8'hba;
frames[8][20][26] = 8'hb6;
frames[8][20][27] = 8'hb6;
frames[8][20][28] = 8'h8d;
frames[8][20][29] = 8'h44;
frames[8][20][30] = 8'hb1;
frames[8][20][31] = 8'hb1;
frames[8][20][32] = 8'hd1;
frames[8][20][33] = 8'hd1;
frames[8][20][34] = 8'hd1;
frames[8][20][35] = 8'hd1;
frames[8][20][36] = 8'hb1;
frames[8][20][37] = 8'hb1;
frames[8][20][38] = 8'hb1;
frames[8][20][39] = 8'hb1;
frames[8][21][0] = 8'hac;
frames[8][21][1] = 8'hac;
frames[8][21][2] = 8'hb1;
frames[8][21][3] = 8'hd1;
frames[8][21][4] = 8'hd1;
frames[8][21][5] = 8'hd1;
frames[8][21][6] = 8'hd5;
frames[8][21][7] = 8'hd5;
frames[8][21][8] = 8'hb1;
frames[8][21][9] = 8'hb1;
frames[8][21][10] = 8'h8d;
frames[8][21][11] = 8'h8d;
frames[8][21][12] = 8'h91;
frames[8][21][13] = 8'h8d;
frames[8][21][14] = 8'h8d;
frames[8][21][15] = 8'h8d;
frames[8][21][16] = 8'ha8;
frames[8][21][17] = 8'h64;
frames[8][21][18] = 8'ha8;
frames[8][21][19] = 8'ha4;
frames[8][21][20] = 8'h8d;
frames[8][21][21] = 8'hb1;
frames[8][21][22] = 8'hb6;
frames[8][21][23] = 8'hb6;
frames[8][21][24] = 8'hb6;
frames[8][21][25] = 8'hb6;
frames[8][21][26] = 8'hb2;
frames[8][21][27] = 8'hb2;
frames[8][21][28] = 8'h91;
frames[8][21][29] = 8'h44;
frames[8][21][30] = 8'had;
frames[8][21][31] = 8'hb1;
frames[8][21][32] = 8'hb1;
frames[8][21][33] = 8'hd1;
frames[8][21][34] = 8'hb1;
frames[8][21][35] = 8'hd1;
frames[8][21][36] = 8'hb1;
frames[8][21][37] = 8'hb1;
frames[8][21][38] = 8'hb1;
frames[8][21][39] = 8'hb1;
frames[8][22][0] = 8'hac;
frames[8][22][1] = 8'hac;
frames[8][22][2] = 8'hb1;
frames[8][22][3] = 8'hd5;
frames[8][22][4] = 8'hd5;
frames[8][22][5] = 8'hd5;
frames[8][22][6] = 8'hd5;
frames[8][22][7] = 8'hd6;
frames[8][22][8] = 8'hd1;
frames[8][22][9] = 8'hb1;
frames[8][22][10] = 8'h91;
frames[8][22][11] = 8'hb1;
frames[8][22][12] = 8'h8d;
frames[8][22][13] = 8'h6d;
frames[8][22][14] = 8'h8d;
frames[8][22][15] = 8'h8d;
frames[8][22][16] = 8'h88;
frames[8][22][17] = 8'h64;
frames[8][22][18] = 8'ha4;
frames[8][22][19] = 8'ha8;
frames[8][22][20] = 8'h8d;
frames[8][22][21] = 8'hb1;
frames[8][22][22] = 8'h91;
frames[8][22][23] = 8'h91;
frames[8][22][24] = 8'h91;
frames[8][22][25] = 8'h91;
frames[8][22][26] = 8'hb1;
frames[8][22][27] = 8'hb1;
frames[8][22][28] = 8'h91;
frames[8][22][29] = 8'h24;
frames[8][22][30] = 8'h8d;
frames[8][22][31] = 8'hb1;
frames[8][22][32] = 8'hb1;
frames[8][22][33] = 8'hb1;
frames[8][22][34] = 8'hb1;
frames[8][22][35] = 8'hd1;
frames[8][22][36] = 8'hb1;
frames[8][22][37] = 8'hb1;
frames[8][22][38] = 8'hb1;
frames[8][22][39] = 8'hb1;
frames[8][23][0] = 8'hac;
frames[8][23][1] = 8'hac;
frames[8][23][2] = 8'hac;
frames[8][23][3] = 8'hb1;
frames[8][23][4] = 8'hb1;
frames[8][23][5] = 8'hb1;
frames[8][23][6] = 8'hd1;
frames[8][23][7] = 8'hd1;
frames[8][23][8] = 8'hb1;
frames[8][23][9] = 8'had;
frames[8][23][10] = 8'h68;
frames[8][23][11] = 8'h8d;
frames[8][23][12] = 8'h8d;
frames[8][23][13] = 8'h8d;
frames[8][23][14] = 8'h8d;
frames[8][23][15] = 8'h8d;
frames[8][23][16] = 8'h89;
frames[8][23][17] = 8'h89;
frames[8][23][18] = 8'h84;
frames[8][23][19] = 8'h84;
frames[8][23][20] = 8'h8d;
frames[8][23][21] = 8'h8d;
frames[8][23][22] = 8'h6d;
frames[8][23][23] = 8'h6d;
frames[8][23][24] = 8'h6d;
frames[8][23][25] = 8'h6d;
frames[8][23][26] = 8'h6d;
frames[8][23][27] = 8'h6d;
frames[8][23][28] = 8'h44;
frames[8][23][29] = 8'h00;
frames[8][23][30] = 8'h8d;
frames[8][23][31] = 8'hb1;
frames[8][23][32] = 8'hd1;
frames[8][23][33] = 8'hb1;
frames[8][23][34] = 8'hb1;
frames[8][23][35] = 8'hd1;
frames[8][23][36] = 8'hb1;
frames[8][23][37] = 8'hb1;
frames[8][23][38] = 8'hb1;
frames[8][23][39] = 8'hb1;
frames[8][24][0] = 8'hac;
frames[8][24][1] = 8'hac;
frames[8][24][2] = 8'hac;
frames[8][24][3] = 8'hac;
frames[8][24][4] = 8'hac;
frames[8][24][5] = 8'hd1;
frames[8][24][6] = 8'hd1;
frames[8][24][7] = 8'hd1;
frames[8][24][8] = 8'hb1;
frames[8][24][9] = 8'hac;
frames[8][24][10] = 8'h20;
frames[8][24][11] = 8'h69;
frames[8][24][12] = 8'h8d;
frames[8][24][13] = 8'h44;
frames[8][24][14] = 8'h44;
frames[8][24][15] = 8'h68;
frames[8][24][16] = 8'h8d;
frames[8][24][17] = 8'h44;
frames[8][24][18] = 8'h44;
frames[8][24][19] = 8'h68;
frames[8][24][20] = 8'h68;
frames[8][24][21] = 8'h69;
frames[8][24][22] = 8'h69;
frames[8][24][23] = 8'h69;
frames[8][24][24] = 8'h69;
frames[8][24][25] = 8'h69;
frames[8][24][26] = 8'h6d;
frames[8][24][27] = 8'h6d;
frames[8][24][28] = 8'h6d;
frames[8][24][29] = 8'h8d;
frames[8][24][30] = 8'hb1;
frames[8][24][31] = 8'hb1;
frames[8][24][32] = 8'hb1;
frames[8][24][33] = 8'hb1;
frames[8][24][34] = 8'hb1;
frames[8][24][35] = 8'hb1;
frames[8][24][36] = 8'hb1;
frames[8][24][37] = 8'hb1;
frames[8][24][38] = 8'hb1;
frames[8][24][39] = 8'hb1;
frames[8][25][0] = 8'hac;
frames[8][25][1] = 8'hac;
frames[8][25][2] = 8'hac;
frames[8][25][3] = 8'hac;
frames[8][25][4] = 8'hb0;
frames[8][25][5] = 8'hb1;
frames[8][25][6] = 8'hd1;
frames[8][25][7] = 8'hd1;
frames[8][25][8] = 8'hd1;
frames[8][25][9] = 8'hd1;
frames[8][25][10] = 8'h8d;
frames[8][25][11] = 8'hb1;
frames[8][25][12] = 8'h8d;
frames[8][25][13] = 8'h8d;
frames[8][25][14] = 8'h8d;
frames[8][25][15] = 8'h8d;
frames[8][25][16] = 8'hb6;
frames[8][25][17] = 8'hb1;
frames[8][25][18] = 8'hb1;
frames[8][25][19] = 8'hb1;
frames[8][25][20] = 8'hb1;
frames[8][25][21] = 8'hb1;
frames[8][25][22] = 8'hd5;
frames[8][25][23] = 8'hd5;
frames[8][25][24] = 8'hd1;
frames[8][25][25] = 8'hd1;
frames[8][25][26] = 8'hd1;
frames[8][25][27] = 8'hd1;
frames[8][25][28] = 8'hd1;
frames[8][25][29] = 8'hd1;
frames[8][25][30] = 8'hb1;
frames[8][25][31] = 8'hb1;
frames[8][25][32] = 8'hb1;
frames[8][25][33] = 8'hb1;
frames[8][25][34] = 8'hb1;
frames[8][25][35] = 8'hb1;
frames[8][25][36] = 8'hb1;
frames[8][25][37] = 8'hb1;
frames[8][25][38] = 8'hb1;
frames[8][25][39] = 8'hb1;
frames[8][26][0] = 8'h8c;
frames[8][26][1] = 8'hac;
frames[8][26][2] = 8'hac;
frames[8][26][3] = 8'hac;
frames[8][26][4] = 8'hac;
frames[8][26][5] = 8'hb1;
frames[8][26][6] = 8'hd1;
frames[8][26][7] = 8'hd1;
frames[8][26][8] = 8'hd1;
frames[8][26][9] = 8'hd1;
frames[8][26][10] = 8'hb1;
frames[8][26][11] = 8'hac;
frames[8][26][12] = 8'hac;
frames[8][26][13] = 8'hb1;
frames[8][26][14] = 8'hb1;
frames[8][26][15] = 8'hb1;
frames[8][26][16] = 8'hb1;
frames[8][26][17] = 8'hb1;
frames[8][26][18] = 8'hb1;
frames[8][26][19] = 8'hd6;
frames[8][26][20] = 8'hd6;
frames[8][26][21] = 8'hd6;
frames[8][26][22] = 8'hd6;
frames[8][26][23] = 8'hd6;
frames[8][26][24] = 8'hd1;
frames[8][26][25] = 8'hd1;
frames[8][26][26] = 8'hd1;
frames[8][26][27] = 8'hb1;
frames[8][26][28] = 8'hb1;
frames[8][26][29] = 8'hb1;
frames[8][26][30] = 8'hb1;
frames[8][26][31] = 8'hb1;
frames[8][26][32] = 8'hb1;
frames[8][26][33] = 8'hb1;
frames[8][26][34] = 8'hb1;
frames[8][26][35] = 8'hb1;
frames[8][26][36] = 8'hb1;
frames[8][26][37] = 8'hb1;
frames[8][26][38] = 8'hb1;
frames[8][26][39] = 8'hb1;
frames[8][27][0] = 8'h8c;
frames[8][27][1] = 8'h8c;
frames[8][27][2] = 8'hac;
frames[8][27][3] = 8'hac;
frames[8][27][4] = 8'hac;
frames[8][27][5] = 8'hb1;
frames[8][27][6] = 8'hd1;
frames[8][27][7] = 8'hd1;
frames[8][27][8] = 8'hd1;
frames[8][27][9] = 8'hd1;
frames[8][27][10] = 8'hd1;
frames[8][27][11] = 8'hb1;
frames[8][27][12] = 8'hb1;
frames[8][27][13] = 8'hb1;
frames[8][27][14] = 8'hb1;
frames[8][27][15] = 8'hb1;
frames[8][27][16] = 8'hac;
frames[8][27][17] = 8'hac;
frames[8][27][18] = 8'hb1;
frames[8][27][19] = 8'hd5;
frames[8][27][20] = 8'hd6;
frames[8][27][21] = 8'hd6;
frames[8][27][22] = 8'hda;
frames[8][27][23] = 8'hd6;
frames[8][27][24] = 8'hd1;
frames[8][27][25] = 8'hb1;
frames[8][27][26] = 8'hb1;
frames[8][27][27] = 8'hb1;
frames[8][27][28] = 8'hb1;
frames[8][27][29] = 8'hb1;
frames[8][27][30] = 8'hb1;
frames[8][27][31] = 8'hb1;
frames[8][27][32] = 8'hb1;
frames[8][27][33] = 8'hb1;
frames[8][27][34] = 8'hb1;
frames[8][27][35] = 8'hb1;
frames[8][27][36] = 8'hb1;
frames[8][27][37] = 8'hb1;
frames[8][27][38] = 8'hb1;
frames[8][27][39] = 8'hb1;
frames[8][28][0] = 8'h88;
frames[8][28][1] = 8'h8c;
frames[8][28][2] = 8'h8c;
frames[8][28][3] = 8'h8c;
frames[8][28][4] = 8'hac;
frames[8][28][5] = 8'hac;
frames[8][28][6] = 8'hb1;
frames[8][28][7] = 8'hb1;
frames[8][28][8] = 8'hd1;
frames[8][28][9] = 8'hd1;
frames[8][28][10] = 8'hb1;
frames[8][28][11] = 8'hb1;
frames[8][28][12] = 8'hb1;
frames[8][28][13] = 8'hb1;
frames[8][28][14] = 8'hb1;
frames[8][28][15] = 8'hb1;
frames[8][28][16] = 8'hac;
frames[8][28][17] = 8'h8c;
frames[8][28][18] = 8'hac;
frames[8][28][19] = 8'had;
frames[8][28][20] = 8'had;
frames[8][28][21] = 8'hb1;
frames[8][28][22] = 8'hd1;
frames[8][28][23] = 8'hd5;
frames[8][28][24] = 8'hb1;
frames[8][28][25] = 8'hb1;
frames[8][28][26] = 8'hb1;
frames[8][28][27] = 8'hb1;
frames[8][28][28] = 8'hb1;
frames[8][28][29] = 8'hb1;
frames[8][28][30] = 8'hb1;
frames[8][28][31] = 8'hb1;
frames[8][28][32] = 8'hb1;
frames[8][28][33] = 8'hb1;
frames[8][28][34] = 8'hb1;
frames[8][28][35] = 8'hb1;
frames[8][28][36] = 8'hb1;
frames[8][28][37] = 8'hb1;
frames[8][28][38] = 8'hb1;
frames[8][28][39] = 8'had;
frames[8][29][0] = 8'h88;
frames[8][29][1] = 8'h8c;
frames[8][29][2] = 8'h8c;
frames[8][29][3] = 8'h8c;
frames[8][29][4] = 8'hac;
frames[8][29][5] = 8'hac;
frames[8][29][6] = 8'hac;
frames[8][29][7] = 8'hb1;
frames[8][29][8] = 8'hd1;
frames[8][29][9] = 8'hb1;
frames[8][29][10] = 8'hb1;
frames[8][29][11] = 8'hb1;
frames[8][29][12] = 8'had;
frames[8][29][13] = 8'hb1;
frames[8][29][14] = 8'hb1;
frames[8][29][15] = 8'hb1;
frames[8][29][16] = 8'hac;
frames[8][29][17] = 8'h8c;
frames[8][29][18] = 8'h8c;
frames[8][29][19] = 8'h8c;
frames[8][29][20] = 8'h8c;
frames[8][29][21] = 8'h8c;
frames[8][29][22] = 8'had;
frames[8][29][23] = 8'hb1;
frames[8][29][24] = 8'hb1;
frames[8][29][25] = 8'hb1;
frames[8][29][26] = 8'hb1;
frames[8][29][27] = 8'hb1;
frames[8][29][28] = 8'hb1;
frames[8][29][29] = 8'hb1;
frames[8][29][30] = 8'hb1;
frames[8][29][31] = 8'hb1;
frames[8][29][32] = 8'hb1;
frames[8][29][33] = 8'hb1;
frames[8][29][34] = 8'hb1;
frames[8][29][35] = 8'hb1;
frames[8][29][36] = 8'hb1;
frames[8][29][37] = 8'hb1;
frames[8][29][38] = 8'hb1;
frames[8][29][39] = 8'hb1;
frames[9][0][0] = 8'hd6;
frames[9][0][1] = 8'hd6;
frames[9][0][2] = 8'hd6;
frames[9][0][3] = 8'hd6;
frames[9][0][4] = 8'hb6;
frames[9][0][5] = 8'h24;
frames[9][0][6] = 8'h00;
frames[9][0][7] = 8'h00;
frames[9][0][8] = 8'h00;
frames[9][0][9] = 8'h00;
frames[9][0][10] = 8'h00;
frames[9][0][11] = 8'h00;
frames[9][0][12] = 8'h00;
frames[9][0][13] = 8'h00;
frames[9][0][14] = 8'h00;
frames[9][0][15] = 8'h00;
frames[9][0][16] = 8'h44;
frames[9][0][17] = 8'h69;
frames[9][0][18] = 8'had;
frames[9][0][19] = 8'had;
frames[9][0][20] = 8'had;
frames[9][0][21] = 8'had;
frames[9][0][22] = 8'had;
frames[9][0][23] = 8'had;
frames[9][0][24] = 8'had;
frames[9][0][25] = 8'had;
frames[9][0][26] = 8'h8d;
frames[9][0][27] = 8'h64;
frames[9][0][28] = 8'h68;
frames[9][0][29] = 8'had;
frames[9][0][30] = 8'hd2;
frames[9][0][31] = 8'hd6;
frames[9][0][32] = 8'hd6;
frames[9][0][33] = 8'hd6;
frames[9][0][34] = 8'hb2;
frames[9][0][35] = 8'hd6;
frames[9][0][36] = 8'hd6;
frames[9][0][37] = 8'hb6;
frames[9][0][38] = 8'hd6;
frames[9][0][39] = 8'hd6;
frames[9][1][0] = 8'hb6;
frames[9][1][1] = 8'hd6;
frames[9][1][2] = 8'hb6;
frames[9][1][3] = 8'hb6;
frames[9][1][4] = 8'h92;
frames[9][1][5] = 8'h00;
frames[9][1][6] = 8'h00;
frames[9][1][7] = 8'h00;
frames[9][1][8] = 8'h00;
frames[9][1][9] = 8'h00;
frames[9][1][10] = 8'h00;
frames[9][1][11] = 8'h00;
frames[9][1][12] = 8'h00;
frames[9][1][13] = 8'h00;
frames[9][1][14] = 8'h00;
frames[9][1][15] = 8'h00;
frames[9][1][16] = 8'h00;
frames[9][1][17] = 8'h00;
frames[9][1][18] = 8'h20;
frames[9][1][19] = 8'h44;
frames[9][1][20] = 8'h89;
frames[9][1][21] = 8'had;
frames[9][1][22] = 8'had;
frames[9][1][23] = 8'had;
frames[9][1][24] = 8'had;
frames[9][1][25] = 8'had;
frames[9][1][26] = 8'had;
frames[9][1][27] = 8'had;
frames[9][1][28] = 8'h89;
frames[9][1][29] = 8'had;
frames[9][1][30] = 8'hb2;
frames[9][1][31] = 8'hd6;
frames[9][1][32] = 8'hd6;
frames[9][1][33] = 8'hd6;
frames[9][1][34] = 8'hb2;
frames[9][1][35] = 8'hd6;
frames[9][1][36] = 8'hdb;
frames[9][1][37] = 8'hda;
frames[9][1][38] = 8'hda;
frames[9][1][39] = 8'hdb;
frames[9][2][0] = 8'hb6;
frames[9][2][1] = 8'hb6;
frames[9][2][2] = 8'hb6;
frames[9][2][3] = 8'hb6;
frames[9][2][4] = 8'h6d;
frames[9][2][5] = 8'h00;
frames[9][2][6] = 8'h00;
frames[9][2][7] = 8'h00;
frames[9][2][8] = 8'h00;
frames[9][2][9] = 8'h00;
frames[9][2][10] = 8'h00;
frames[9][2][11] = 8'h00;
frames[9][2][12] = 8'h00;
frames[9][2][13] = 8'h00;
frames[9][2][14] = 8'h00;
frames[9][2][15] = 8'h00;
frames[9][2][16] = 8'h00;
frames[9][2][17] = 8'h00;
frames[9][2][18] = 8'h00;
frames[9][2][19] = 8'h00;
frames[9][2][20] = 8'h00;
frames[9][2][21] = 8'h20;
frames[9][2][22] = 8'h68;
frames[9][2][23] = 8'had;
frames[9][2][24] = 8'had;
frames[9][2][25] = 8'had;
frames[9][2][26] = 8'had;
frames[9][2][27] = 8'had;
frames[9][2][28] = 8'hd1;
frames[9][2][29] = 8'had;
frames[9][2][30] = 8'hb2;
frames[9][2][31] = 8'hd6;
frames[9][2][32] = 8'hd6;
frames[9][2][33] = 8'hd6;
frames[9][2][34] = 8'hb2;
frames[9][2][35] = 8'hd6;
frames[9][2][36] = 8'hfb;
frames[9][2][37] = 8'h92;
frames[9][2][38] = 8'hb2;
frames[9][2][39] = 8'hdb;
frames[9][3][0] = 8'hb2;
frames[9][3][1] = 8'hb6;
frames[9][3][2] = 8'hb6;
frames[9][3][3] = 8'hb6;
frames[9][3][4] = 8'h69;
frames[9][3][5] = 8'h00;
frames[9][3][6] = 8'h00;
frames[9][3][7] = 8'h00;
frames[9][3][8] = 8'h00;
frames[9][3][9] = 8'h00;
frames[9][3][10] = 8'h00;
frames[9][3][11] = 8'h00;
frames[9][3][12] = 8'h00;
frames[9][3][13] = 8'h00;
frames[9][3][14] = 8'h00;
frames[9][3][15] = 8'h00;
frames[9][3][16] = 8'h00;
frames[9][3][17] = 8'h00;
frames[9][3][18] = 8'h00;
frames[9][3][19] = 8'h00;
frames[9][3][20] = 8'h00;
frames[9][3][21] = 8'h00;
frames[9][3][22] = 8'h20;
frames[9][3][23] = 8'h8d;
frames[9][3][24] = 8'had;
frames[9][3][25] = 8'had;
frames[9][3][26] = 8'had;
frames[9][3][27] = 8'had;
frames[9][3][28] = 8'hd1;
frames[9][3][29] = 8'hcd;
frames[9][3][30] = 8'hb2;
frames[9][3][31] = 8'hd6;
frames[9][3][32] = 8'hd6;
frames[9][3][33] = 8'hd6;
frames[9][3][34] = 8'hb2;
frames[9][3][35] = 8'hd6;
frames[9][3][36] = 8'hdb;
frames[9][3][37] = 8'hb2;
frames[9][3][38] = 8'hd6;
frames[9][3][39] = 8'hfb;
frames[9][4][0] = 8'hb2;
frames[9][4][1] = 8'hb6;
frames[9][4][2] = 8'hb6;
frames[9][4][3] = 8'hb6;
frames[9][4][4] = 8'h49;
frames[9][4][5] = 8'h00;
frames[9][4][6] = 8'h00;
frames[9][4][7] = 8'h00;
frames[9][4][8] = 8'h00;
frames[9][4][9] = 8'h00;
frames[9][4][10] = 8'h00;
frames[9][4][11] = 8'h00;
frames[9][4][12] = 8'h00;
frames[9][4][13] = 8'h00;
frames[9][4][14] = 8'h00;
frames[9][4][15] = 8'h00;
frames[9][4][16] = 8'h00;
frames[9][4][17] = 8'h00;
frames[9][4][18] = 8'h00;
frames[9][4][19] = 8'h00;
frames[9][4][20] = 8'h00;
frames[9][4][21] = 8'h00;
frames[9][4][22] = 8'h00;
frames[9][4][23] = 8'h44;
frames[9][4][24] = 8'hb1;
frames[9][4][25] = 8'had;
frames[9][4][26] = 8'had;
frames[9][4][27] = 8'had;
frames[9][4][28] = 8'had;
frames[9][4][29] = 8'had;
frames[9][4][30] = 8'hb2;
frames[9][4][31] = 8'hd6;
frames[9][4][32] = 8'hd6;
frames[9][4][33] = 8'hd6;
frames[9][4][34] = 8'hb2;
frames[9][4][35] = 8'hd6;
frames[9][4][36] = 8'hfb;
frames[9][4][37] = 8'hb6;
frames[9][4][38] = 8'hda;
frames[9][4][39] = 8'hdb;
frames[9][5][0] = 8'hb2;
frames[9][5][1] = 8'hb6;
frames[9][5][2] = 8'hb6;
frames[9][5][3] = 8'hb6;
frames[9][5][4] = 8'h24;
frames[9][5][5] = 8'h00;
frames[9][5][6] = 8'h00;
frames[9][5][7] = 8'h00;
frames[9][5][8] = 8'h00;
frames[9][5][9] = 8'h00;
frames[9][5][10] = 8'h00;
frames[9][5][11] = 8'h00;
frames[9][5][12] = 8'h00;
frames[9][5][13] = 8'h00;
frames[9][5][14] = 8'h00;
frames[9][5][15] = 8'h00;
frames[9][5][16] = 8'h00;
frames[9][5][17] = 8'h00;
frames[9][5][18] = 8'h00;
frames[9][5][19] = 8'h00;
frames[9][5][20] = 8'h00;
frames[9][5][21] = 8'h00;
frames[9][5][22] = 8'h00;
frames[9][5][23] = 8'h00;
frames[9][5][24] = 8'h68;
frames[9][5][25] = 8'had;
frames[9][5][26] = 8'had;
frames[9][5][27] = 8'had;
frames[9][5][28] = 8'had;
frames[9][5][29] = 8'had;
frames[9][5][30] = 8'hb1;
frames[9][5][31] = 8'hd6;
frames[9][5][32] = 8'hd6;
frames[9][5][33] = 8'hd6;
frames[9][5][34] = 8'hb2;
frames[9][5][35] = 8'hd6;
frames[9][5][36] = 8'hd6;
frames[9][5][37] = 8'hda;
frames[9][5][38] = 8'hdb;
frames[9][5][39] = 8'hd6;
frames[9][6][0] = 8'h92;
frames[9][6][1] = 8'hb2;
frames[9][6][2] = 8'h92;
frames[9][6][3] = 8'h92;
frames[9][6][4] = 8'h49;
frames[9][6][5] = 8'h00;
frames[9][6][6] = 8'h00;
frames[9][6][7] = 8'h00;
frames[9][6][8] = 8'h00;
frames[9][6][9] = 8'h00;
frames[9][6][10] = 8'h00;
frames[9][6][11] = 8'h00;
frames[9][6][12] = 8'h00;
frames[9][6][13] = 8'h00;
frames[9][6][14] = 8'h00;
frames[9][6][15] = 8'h00;
frames[9][6][16] = 8'h00;
frames[9][6][17] = 8'h00;
frames[9][6][18] = 8'h00;
frames[9][6][19] = 8'h00;
frames[9][6][20] = 8'h00;
frames[9][6][21] = 8'h00;
frames[9][6][22] = 8'h00;
frames[9][6][23] = 8'h00;
frames[9][6][24] = 8'h44;
frames[9][6][25] = 8'h8d;
frames[9][6][26] = 8'had;
frames[9][6][27] = 8'had;
frames[9][6][28] = 8'had;
frames[9][6][29] = 8'had;
frames[9][6][30] = 8'hb1;
frames[9][6][31] = 8'hd6;
frames[9][6][32] = 8'hd6;
frames[9][6][33] = 8'hd6;
frames[9][6][34] = 8'hb2;
frames[9][6][35] = 8'hd6;
frames[9][6][36] = 8'hd6;
frames[9][6][37] = 8'h91;
frames[9][6][38] = 8'hd6;
frames[9][6][39] = 8'hd6;
frames[9][7][0] = 8'h71;
frames[9][7][1] = 8'h71;
frames[9][7][2] = 8'h71;
frames[9][7][3] = 8'h72;
frames[9][7][4] = 8'h92;
frames[9][7][5] = 8'h92;
frames[9][7][6] = 8'h91;
frames[9][7][7] = 8'h49;
frames[9][7][8] = 8'h00;
frames[9][7][9] = 8'h00;
frames[9][7][10] = 8'h00;
frames[9][7][11] = 8'h00;
frames[9][7][12] = 8'h00;
frames[9][7][13] = 8'h00;
frames[9][7][14] = 8'h00;
frames[9][7][15] = 8'h00;
frames[9][7][16] = 8'h00;
frames[9][7][17] = 8'h00;
frames[9][7][18] = 8'h00;
frames[9][7][19] = 8'h00;
frames[9][7][20] = 8'h00;
frames[9][7][21] = 8'h00;
frames[9][7][22] = 8'h00;
frames[9][7][23] = 8'h00;
frames[9][7][24] = 8'h44;
frames[9][7][25] = 8'h64;
frames[9][7][26] = 8'h89;
frames[9][7][27] = 8'had;
frames[9][7][28] = 8'had;
frames[9][7][29] = 8'had;
frames[9][7][30] = 8'h8d;
frames[9][7][31] = 8'hd2;
frames[9][7][32] = 8'hd6;
frames[9][7][33] = 8'hd6;
frames[9][7][34] = 8'hb2;
frames[9][7][35] = 8'hd6;
frames[9][7][36] = 8'hd6;
frames[9][7][37] = 8'h91;
frames[9][7][38] = 8'hd6;
frames[9][7][39] = 8'hd6;
frames[9][8][0] = 8'h91;
frames[9][8][1] = 8'h92;
frames[9][8][2] = 8'hb6;
frames[9][8][3] = 8'hb6;
frames[9][8][4] = 8'hd6;
frames[9][8][5] = 8'hd6;
frames[9][8][6] = 8'hda;
frames[9][8][7] = 8'hda;
frames[9][8][8] = 8'h92;
frames[9][8][9] = 8'h44;
frames[9][8][10] = 8'h20;
frames[9][8][11] = 8'h20;
frames[9][8][12] = 8'h20;
frames[9][8][13] = 8'h20;
frames[9][8][14] = 8'h20;
frames[9][8][15] = 8'h24;
frames[9][8][16] = 8'h24;
frames[9][8][17] = 8'h24;
frames[9][8][18] = 8'h24;
frames[9][8][19] = 8'h48;
frames[9][8][20] = 8'h48;
frames[9][8][21] = 8'h48;
frames[9][8][22] = 8'h48;
frames[9][8][23] = 8'h48;
frames[9][8][24] = 8'h44;
frames[9][8][25] = 8'h44;
frames[9][8][26] = 8'h88;
frames[9][8][27] = 8'had;
frames[9][8][28] = 8'had;
frames[9][8][29] = 8'ha9;
frames[9][8][30] = 8'h69;
frames[9][8][31] = 8'h68;
frames[9][8][32] = 8'h6d;
frames[9][8][33] = 8'h6d;
frames[9][8][34] = 8'h6d;
frames[9][8][35] = 8'h91;
frames[9][8][36] = 8'hd6;
frames[9][8][37] = 8'hda;
frames[9][8][38] = 8'hfa;
frames[9][8][39] = 8'hfb;
frames[9][9][0] = 8'hd6;
frames[9][9][1] = 8'hd6;
frames[9][9][2] = 8'hd6;
frames[9][9][3] = 8'hd6;
frames[9][9][4] = 8'hd6;
frames[9][9][5] = 8'hd6;
frames[9][9][6] = 8'hd6;
frames[9][9][7] = 8'hd6;
frames[9][9][8] = 8'hb6;
frames[9][9][9] = 8'h91;
frames[9][9][10] = 8'h68;
frames[9][9][11] = 8'h64;
frames[9][9][12] = 8'h68;
frames[9][9][13] = 8'h88;
frames[9][9][14] = 8'h68;
frames[9][9][15] = 8'h68;
frames[9][9][16] = 8'h44;
frames[9][9][17] = 8'h44;
frames[9][9][18] = 8'h24;
frames[9][9][19] = 8'h49;
frames[9][9][20] = 8'h49;
frames[9][9][21] = 8'h49;
frames[9][9][22] = 8'h49;
frames[9][9][23] = 8'h69;
frames[9][9][24] = 8'h69;
frames[9][9][25] = 8'h6d;
frames[9][9][26] = 8'h8d;
frames[9][9][27] = 8'had;
frames[9][9][28] = 8'had;
frames[9][9][29] = 8'had;
frames[9][9][30] = 8'h69;
frames[9][9][31] = 8'h20;
frames[9][9][32] = 8'h44;
frames[9][9][33] = 8'h48;
frames[9][9][34] = 8'h49;
frames[9][9][35] = 8'h49;
frames[9][9][36] = 8'hb2;
frames[9][9][37] = 8'hff;
frames[9][9][38] = 8'hff;
frames[9][9][39] = 8'hff;
frames[9][10][0] = 8'hda;
frames[9][10][1] = 8'hda;
frames[9][10][2] = 8'hda;
frames[9][10][3] = 8'hd6;
frames[9][10][4] = 8'hd6;
frames[9][10][5] = 8'hd6;
frames[9][10][6] = 8'hd6;
frames[9][10][7] = 8'hb1;
frames[9][10][8] = 8'hb2;
frames[9][10][9] = 8'h91;
frames[9][10][10] = 8'h88;
frames[9][10][11] = 8'h68;
frames[9][10][12] = 8'h88;
frames[9][10][13] = 8'h88;
frames[9][10][14] = 8'h68;
frames[9][10][15] = 8'h44;
frames[9][10][16] = 8'h24;
frames[9][10][17] = 8'h44;
frames[9][10][18] = 8'h24;
frames[9][10][19] = 8'h24;
frames[9][10][20] = 8'h24;
frames[9][10][21] = 8'h24;
frames[9][10][22] = 8'h8d;
frames[9][10][23] = 8'hd6;
frames[9][10][24] = 8'hd6;
frames[9][10][25] = 8'hda;
frames[9][10][26] = 8'hf6;
frames[9][10][27] = 8'had;
frames[9][10][28] = 8'had;
frames[9][10][29] = 8'hd1;
frames[9][10][30] = 8'hd6;
frames[9][10][31] = 8'hb1;
frames[9][10][32] = 8'h69;
frames[9][10][33] = 8'h49;
frames[9][10][34] = 8'h49;
frames[9][10][35] = 8'h24;
frames[9][10][36] = 8'h8d;
frames[9][10][37] = 8'hff;
frames[9][10][38] = 8'hff;
frames[9][10][39] = 8'hff;
frames[9][11][0] = 8'hd6;
frames[9][11][1] = 8'hd6;
frames[9][11][2] = 8'hd6;
frames[9][11][3] = 8'hd6;
frames[9][11][4] = 8'hd6;
frames[9][11][5] = 8'hd6;
frames[9][11][6] = 8'hd6;
frames[9][11][7] = 8'hb6;
frames[9][11][8] = 8'h91;
frames[9][11][9] = 8'h6d;
frames[9][11][10] = 8'h68;
frames[9][11][11] = 8'h68;
frames[9][11][12] = 8'h88;
frames[9][11][13] = 8'h88;
frames[9][11][14] = 8'h64;
frames[9][11][15] = 8'h40;
frames[9][11][16] = 8'h24;
frames[9][11][17] = 8'h24;
frames[9][11][18] = 8'h24;
frames[9][11][19] = 8'h24;
frames[9][11][20] = 8'h44;
frames[9][11][21] = 8'h92;
frames[9][11][22] = 8'hd6;
frames[9][11][23] = 8'hd6;
frames[9][11][24] = 8'hd6;
frames[9][11][25] = 8'hd6;
frames[9][11][26] = 8'hb1;
frames[9][11][27] = 8'hd1;
frames[9][11][28] = 8'hb1;
frames[9][11][29] = 8'hf6;
frames[9][11][30] = 8'hda;
frames[9][11][31] = 8'hda;
frames[9][11][32] = 8'hd6;
frames[9][11][33] = 8'hb2;
frames[9][11][34] = 8'h92;
frames[9][11][35] = 8'h6d;
frames[9][11][36] = 8'h69;
frames[9][11][37] = 8'hff;
frames[9][11][38] = 8'hff;
frames[9][11][39] = 8'hff;
frames[9][12][0] = 8'hd6;
frames[9][12][1] = 8'hd6;
frames[9][12][2] = 8'hd6;
frames[9][12][3] = 8'hb6;
frames[9][12][4] = 8'hb6;
frames[9][12][5] = 8'hb1;
frames[9][12][6] = 8'hb1;
frames[9][12][7] = 8'h8d;
frames[9][12][8] = 8'h8d;
frames[9][12][9] = 8'h6d;
frames[9][12][10] = 8'h68;
frames[9][12][11] = 8'h88;
frames[9][12][12] = 8'h88;
frames[9][12][13] = 8'h88;
frames[9][12][14] = 8'h64;
frames[9][12][15] = 8'h44;
frames[9][12][16] = 8'h24;
frames[9][12][17] = 8'h24;
frames[9][12][18] = 8'h24;
frames[9][12][19] = 8'h24;
frames[9][12][20] = 8'h48;
frames[9][12][21] = 8'hb1;
frames[9][12][22] = 8'hb1;
frames[9][12][23] = 8'hb5;
frames[9][12][24] = 8'hb5;
frames[9][12][25] = 8'hd5;
frames[9][12][26] = 8'hb1;
frames[9][12][27] = 8'hd5;
frames[9][12][28] = 8'hb5;
frames[9][12][29] = 8'hd6;
frames[9][12][30] = 8'hda;
frames[9][12][31] = 8'hda;
frames[9][12][32] = 8'hda;
frames[9][12][33] = 8'hd6;
frames[9][12][34] = 8'hb6;
frames[9][12][35] = 8'h92;
frames[9][12][36] = 8'h49;
frames[9][12][37] = 8'hdb;
frames[9][12][38] = 8'hff;
frames[9][12][39] = 8'hff;
frames[9][13][0] = 8'hd6;
frames[9][13][1] = 8'hd6;
frames[9][13][2] = 8'hb6;
frames[9][13][3] = 8'hb2;
frames[9][13][4] = 8'hb1;
frames[9][13][5] = 8'hb1;
frames[9][13][6] = 8'h8d;
frames[9][13][7] = 8'h6d;
frames[9][13][8] = 8'h8d;
frames[9][13][9] = 8'h68;
frames[9][13][10] = 8'h68;
frames[9][13][11] = 8'h88;
frames[9][13][12] = 8'h88;
frames[9][13][13] = 8'h88;
frames[9][13][14] = 8'h64;
frames[9][13][15] = 8'h44;
frames[9][13][16] = 8'h24;
frames[9][13][17] = 8'h20;
frames[9][13][18] = 8'h00;
frames[9][13][19] = 8'h00;
frames[9][13][20] = 8'h44;
frames[9][13][21] = 8'h8d;
frames[9][13][22] = 8'h8d;
frames[9][13][23] = 8'hb1;
frames[9][13][24] = 8'hb5;
frames[9][13][25] = 8'hda;
frames[9][13][26] = 8'hda;
frames[9][13][27] = 8'hfa;
frames[9][13][28] = 8'hda;
frames[9][13][29] = 8'hfa;
frames[9][13][30] = 8'hfa;
frames[9][13][31] = 8'hd6;
frames[9][13][32] = 8'hda;
frames[9][13][33] = 8'hda;
frames[9][13][34] = 8'hd6;
frames[9][13][35] = 8'hb6;
frames[9][13][36] = 8'h49;
frames[9][13][37] = 8'hb6;
frames[9][13][38] = 8'hff;
frames[9][13][39] = 8'hff;
frames[9][14][0] = 8'hd6;
frames[9][14][1] = 8'hb6;
frames[9][14][2] = 8'hb6;
frames[9][14][3] = 8'hb1;
frames[9][14][4] = 8'h91;
frames[9][14][5] = 8'h91;
frames[9][14][6] = 8'h6d;
frames[9][14][7] = 8'h6d;
frames[9][14][8] = 8'hb1;
frames[9][14][9] = 8'h48;
frames[9][14][10] = 8'h68;
frames[9][14][11] = 8'h68;
frames[9][14][12] = 8'h88;
frames[9][14][13] = 8'h68;
frames[9][14][14] = 8'h44;
frames[9][14][15] = 8'h44;
frames[9][14][16] = 8'h24;
frames[9][14][17] = 8'h20;
frames[9][14][18] = 8'h00;
frames[9][14][19] = 8'h00;
frames[9][14][20] = 8'h20;
frames[9][14][21] = 8'h69;
frames[9][14][22] = 8'h91;
frames[9][14][23] = 8'hb5;
frames[9][14][24] = 8'hd5;
frames[9][14][25] = 8'hd5;
frames[9][14][26] = 8'hd6;
frames[9][14][27] = 8'hfa;
frames[9][14][28] = 8'hfa;
frames[9][14][29] = 8'hfa;
frames[9][14][30] = 8'hfa;
frames[9][14][31] = 8'hfa;
frames[9][14][32] = 8'hda;
frames[9][14][33] = 8'hda;
frames[9][14][34] = 8'hb6;
frames[9][14][35] = 8'hb6;
frames[9][14][36] = 8'h49;
frames[9][14][37] = 8'h92;
frames[9][14][38] = 8'hff;
frames[9][14][39] = 8'hff;
frames[9][15][0] = 8'h91;
frames[9][15][1] = 8'h91;
frames[9][15][2] = 8'h91;
frames[9][15][3] = 8'h91;
frames[9][15][4] = 8'h91;
frames[9][15][5] = 8'hb1;
frames[9][15][6] = 8'h8d;
frames[9][15][7] = 8'h8d;
frames[9][15][8] = 8'hb2;
frames[9][15][9] = 8'h44;
frames[9][15][10] = 8'h68;
frames[9][15][11] = 8'h68;
frames[9][15][12] = 8'h8d;
frames[9][15][13] = 8'h68;
frames[9][15][14] = 8'h44;
frames[9][15][15] = 8'h44;
frames[9][15][16] = 8'h24;
frames[9][15][17] = 8'h20;
frames[9][15][18] = 8'h20;
frames[9][15][19] = 8'h24;
frames[9][15][20] = 8'h24;
frames[9][15][21] = 8'h24;
frames[9][15][22] = 8'h68;
frames[9][15][23] = 8'hb1;
frames[9][15][24] = 8'hd6;
frames[9][15][25] = 8'hb5;
frames[9][15][26] = 8'hd6;
frames[9][15][27] = 8'hd6;
frames[9][15][28] = 8'hda;
frames[9][15][29] = 8'hda;
frames[9][15][30] = 8'hd6;
frames[9][15][31] = 8'hfa;
frames[9][15][32] = 8'hda;
frames[9][15][33] = 8'hb1;
frames[9][15][34] = 8'h91;
frames[9][15][35] = 8'hb6;
frames[9][15][36] = 8'h6d;
frames[9][15][37] = 8'h6d;
frames[9][15][38] = 8'hff;
frames[9][15][39] = 8'hff;
frames[9][16][0] = 8'h8d;
frames[9][16][1] = 8'h91;
frames[9][16][2] = 8'h8d;
frames[9][16][3] = 8'h8d;
frames[9][16][4] = 8'h8d;
frames[9][16][5] = 8'hd6;
frames[9][16][6] = 8'hd5;
frames[9][16][7] = 8'hd5;
frames[9][16][8] = 8'hd1;
frames[9][16][9] = 8'h8d;
frames[9][16][10] = 8'h8c;
frames[9][16][11] = 8'h8c;
frames[9][16][12] = 8'h8d;
frames[9][16][13] = 8'h68;
frames[9][16][14] = 8'h44;
frames[9][16][15] = 8'h44;
frames[9][16][16] = 8'h44;
frames[9][16][17] = 8'h24;
frames[9][16][18] = 8'h24;
frames[9][16][19] = 8'h24;
frames[9][16][20] = 8'h24;
frames[9][16][21] = 8'h24;
frames[9][16][22] = 8'h24;
frames[9][16][23] = 8'h44;
frames[9][16][24] = 8'h6d;
frames[9][16][25] = 8'h91;
frames[9][16][26] = 8'hb1;
frames[9][16][27] = 8'hb5;
frames[9][16][28] = 8'hb6;
frames[9][16][29] = 8'hb6;
frames[9][16][30] = 8'hb6;
frames[9][16][31] = 8'h91;
frames[9][16][32] = 8'h6d;
frames[9][16][33] = 8'h6d;
frames[9][16][34] = 8'h92;
frames[9][16][35] = 8'hb6;
frames[9][16][36] = 8'h6d;
frames[9][16][37] = 8'h6d;
frames[9][16][38] = 8'hff;
frames[9][16][39] = 8'hff;
frames[9][17][0] = 8'h69;
frames[9][17][1] = 8'h8d;
frames[9][17][2] = 8'h8d;
frames[9][17][3] = 8'hd5;
frames[9][17][4] = 8'hd5;
frames[9][17][5] = 8'hd5;
frames[9][17][6] = 8'hd6;
frames[9][17][7] = 8'hd5;
frames[9][17][8] = 8'hd6;
frames[9][17][9] = 8'hd6;
frames[9][17][10] = 8'hd5;
frames[9][17][11] = 8'hb1;
frames[9][17][12] = 8'h8d;
frames[9][17][13] = 8'h68;
frames[9][17][14] = 8'h44;
frames[9][17][15] = 8'h44;
frames[9][17][16] = 8'h44;
frames[9][17][17] = 8'h44;
frames[9][17][18] = 8'h24;
frames[9][17][19] = 8'h24;
frames[9][17][20] = 8'h24;
frames[9][17][21] = 8'h44;
frames[9][17][22] = 8'h44;
frames[9][17][23] = 8'h44;
frames[9][17][24] = 8'h44;
frames[9][17][25] = 8'h24;
frames[9][17][26] = 8'h44;
frames[9][17][27] = 8'h44;
frames[9][17][28] = 8'h48;
frames[9][17][29] = 8'h44;
frames[9][17][30] = 8'h44;
frames[9][17][31] = 8'h49;
frames[9][17][32] = 8'h6d;
frames[9][17][33] = 8'h92;
frames[9][17][34] = 8'h96;
frames[9][17][35] = 8'hb6;
frames[9][17][36] = 8'h92;
frames[9][17][37] = 8'h49;
frames[9][17][38] = 8'hdb;
frames[9][17][39] = 8'hff;
frames[9][18][0] = 8'h68;
frames[9][18][1] = 8'hb1;
frames[9][18][2] = 8'hd5;
frames[9][18][3] = 8'hd6;
frames[9][18][4] = 8'hd6;
frames[9][18][5] = 8'hd5;
frames[9][18][6] = 8'hd5;
frames[9][18][7] = 8'hd5;
frames[9][18][8] = 8'hd5;
frames[9][18][9] = 8'hd5;
frames[9][18][10] = 8'hd5;
frames[9][18][11] = 8'hb1;
frames[9][18][12] = 8'h8d;
frames[9][18][13] = 8'h68;
frames[9][18][14] = 8'h44;
frames[9][18][15] = 8'h44;
frames[9][18][16] = 8'h44;
frames[9][18][17] = 8'h44;
frames[9][18][18] = 8'h24;
frames[9][18][19] = 8'h24;
frames[9][18][20] = 8'h24;
frames[9][18][21] = 8'h44;
frames[9][18][22] = 8'h44;
frames[9][18][23] = 8'h48;
frames[9][18][24] = 8'h6d;
frames[9][18][25] = 8'h8d;
frames[9][18][26] = 8'hb1;
frames[9][18][27] = 8'hb6;
frames[9][18][28] = 8'hd6;
frames[9][18][29] = 8'hb6;
frames[9][18][30] = 8'hb6;
frames[9][18][31] = 8'hb6;
frames[9][18][32] = 8'hb6;
frames[9][18][33] = 8'hb6;
frames[9][18][34] = 8'h92;
frames[9][18][35] = 8'hb6;
frames[9][18][36] = 8'h92;
frames[9][18][37] = 8'h49;
frames[9][18][38] = 8'hb6;
frames[9][18][39] = 8'hff;
frames[9][19][0] = 8'h88;
frames[9][19][1] = 8'had;
frames[9][19][2] = 8'hd6;
frames[9][19][3] = 8'hda;
frames[9][19][4] = 8'hd6;
frames[9][19][5] = 8'hda;
frames[9][19][6] = 8'hd5;
frames[9][19][7] = 8'hd5;
frames[9][19][8] = 8'hb1;
frames[9][19][9] = 8'hd5;
frames[9][19][10] = 8'hb5;
frames[9][19][11] = 8'hb1;
frames[9][19][12] = 8'h8c;
frames[9][19][13] = 8'h68;
frames[9][19][14] = 8'h64;
frames[9][19][15] = 8'h44;
frames[9][19][16] = 8'h44;
frames[9][19][17] = 8'h44;
frames[9][19][18] = 8'h24;
frames[9][19][19] = 8'h44;
frames[9][19][20] = 8'h44;
frames[9][19][21] = 8'h44;
frames[9][19][22] = 8'h68;
frames[9][19][23] = 8'hb2;
frames[9][19][24] = 8'hd6;
frames[9][19][25] = 8'hd6;
frames[9][19][26] = 8'hd6;
frames[9][19][27] = 8'hd6;
frames[9][19][28] = 8'hd6;
frames[9][19][29] = 8'hd6;
frames[9][19][30] = 8'hda;
frames[9][19][31] = 8'hda;
frames[9][19][32] = 8'hda;
frames[9][19][33] = 8'hd6;
frames[9][19][34] = 8'hb6;
frames[9][19][35] = 8'hb6;
frames[9][19][36] = 8'hb2;
frames[9][19][37] = 8'h49;
frames[9][19][38] = 8'h92;
frames[9][19][39] = 8'hff;
frames[9][20][0] = 8'had;
frames[9][20][1] = 8'hb1;
frames[9][20][2] = 8'hb5;
frames[9][20][3] = 8'hd5;
frames[9][20][4] = 8'hd6;
frames[9][20][5] = 8'hd6;
frames[9][20][6] = 8'hd6;
frames[9][20][7] = 8'hd6;
frames[9][20][8] = 8'hd5;
frames[9][20][9] = 8'hb5;
frames[9][20][10] = 8'hb1;
frames[9][20][11] = 8'hb1;
frames[9][20][12] = 8'h8c;
frames[9][20][13] = 8'h88;
frames[9][20][14] = 8'h64;
frames[9][20][15] = 8'h64;
frames[9][20][16] = 8'h44;
frames[9][20][17] = 8'h44;
frames[9][20][18] = 8'h24;
frames[9][20][19] = 8'h44;
frames[9][20][20] = 8'h44;
frames[9][20][21] = 8'h44;
frames[9][20][22] = 8'hb1;
frames[9][20][23] = 8'hd6;
frames[9][20][24] = 8'hd6;
frames[9][20][25] = 8'hd6;
frames[9][20][26] = 8'hd6;
frames[9][20][27] = 8'hd6;
frames[9][20][28] = 8'hd6;
frames[9][20][29] = 8'hd6;
frames[9][20][30] = 8'hda;
frames[9][20][31] = 8'hda;
frames[9][20][32] = 8'hda;
frames[9][20][33] = 8'hd6;
frames[9][20][34] = 8'hd6;
frames[9][20][35] = 8'hb6;
frames[9][20][36] = 8'hb6;
frames[9][20][37] = 8'h6d;
frames[9][20][38] = 8'h6d;
frames[9][20][39] = 8'hff;
frames[9][21][0] = 8'hb1;
frames[9][21][1] = 8'hb1;
frames[9][21][2] = 8'hd5;
frames[9][21][3] = 8'hfa;
frames[9][21][4] = 8'hda;
frames[9][21][5] = 8'hfa;
frames[9][21][6] = 8'hfa;
frames[9][21][7] = 8'hfa;
frames[9][21][8] = 8'hd6;
frames[9][21][9] = 8'hd5;
frames[9][21][10] = 8'hd5;
frames[9][21][11] = 8'hb1;
frames[9][21][12] = 8'hac;
frames[9][21][13] = 8'h88;
frames[9][21][14] = 8'h68;
frames[9][21][15] = 8'h64;
frames[9][21][16] = 8'h44;
frames[9][21][17] = 8'h44;
frames[9][21][18] = 8'h24;
frames[9][21][19] = 8'h44;
frames[9][21][20] = 8'h44;
frames[9][21][21] = 8'h69;
frames[9][21][22] = 8'hd6;
frames[9][21][23] = 8'hd6;
frames[9][21][24] = 8'hd6;
frames[9][21][25] = 8'hd6;
frames[9][21][26] = 8'hd6;
frames[9][21][27] = 8'hd6;
frames[9][21][28] = 8'hd6;
frames[9][21][29] = 8'hd6;
frames[9][21][30] = 8'hda;
frames[9][21][31] = 8'hda;
frames[9][21][32] = 8'hda;
frames[9][21][33] = 8'hda;
frames[9][21][34] = 8'hd6;
frames[9][21][35] = 8'hd6;
frames[9][21][36] = 8'hb6;
frames[9][21][37] = 8'h6d;
frames[9][21][38] = 8'h49;
frames[9][21][39] = 8'hfb;
frames[9][22][0] = 8'hb2;
frames[9][22][1] = 8'hb2;
frames[9][22][2] = 8'hb1;
frames[9][22][3] = 8'hd6;
frames[9][22][4] = 8'hfa;
frames[9][22][5] = 8'hfa;
frames[9][22][6] = 8'hda;
frames[9][22][7] = 8'hfa;
frames[9][22][8] = 8'hd6;
frames[9][22][9] = 8'hb5;
frames[9][22][10] = 8'hb1;
frames[9][22][11] = 8'hac;
frames[9][22][12] = 8'hac;
frames[9][22][13] = 8'h88;
frames[9][22][14] = 8'h88;
frames[9][22][15] = 8'h64;
frames[9][22][16] = 8'h44;
frames[9][22][17] = 8'h24;
frames[9][22][18] = 8'h24;
frames[9][22][19] = 8'h44;
frames[9][22][20] = 8'h44;
frames[9][22][21] = 8'h69;
frames[9][22][22] = 8'hd6;
frames[9][22][23] = 8'hd6;
frames[9][22][24] = 8'hd6;
frames[9][22][25] = 8'hd6;
frames[9][22][26] = 8'hd6;
frames[9][22][27] = 8'hd6;
frames[9][22][28] = 8'hd6;
frames[9][22][29] = 8'hd6;
frames[9][22][30] = 8'hd6;
frames[9][22][31] = 8'hda;
frames[9][22][32] = 8'hda;
frames[9][22][33] = 8'hda;
frames[9][22][34] = 8'hda;
frames[9][22][35] = 8'hd6;
frames[9][22][36] = 8'hb6;
frames[9][22][37] = 8'h71;
frames[9][22][38] = 8'h48;
frames[9][22][39] = 8'hda;
frames[9][23][0] = 8'hb2;
frames[9][23][1] = 8'hb2;
frames[9][23][2] = 8'hb1;
frames[9][23][3] = 8'h8d;
frames[9][23][4] = 8'hb1;
frames[9][23][5] = 8'hd5;
frames[9][23][6] = 8'hd5;
frames[9][23][7] = 8'hd5;
frames[9][23][8] = 8'hb1;
frames[9][23][9] = 8'had;
frames[9][23][10] = 8'hac;
frames[9][23][11] = 8'hac;
frames[9][23][12] = 8'hac;
frames[9][23][13] = 8'h88;
frames[9][23][14] = 8'h68;
frames[9][23][15] = 8'h64;
frames[9][23][16] = 8'h44;
frames[9][23][17] = 8'h24;
frames[9][23][18] = 8'h44;
frames[9][23][19] = 8'h44;
frames[9][23][20] = 8'h44;
frames[9][23][21] = 8'h44;
frames[9][23][22] = 8'hb1;
frames[9][23][23] = 8'hd6;
frames[9][23][24] = 8'hd6;
frames[9][23][25] = 8'hd6;
frames[9][23][26] = 8'hd6;
frames[9][23][27] = 8'hd6;
frames[9][23][28] = 8'hd6;
frames[9][23][29] = 8'hd6;
frames[9][23][30] = 8'hd6;
frames[9][23][31] = 8'hda;
frames[9][23][32] = 8'hda;
frames[9][23][33] = 8'hda;
frames[9][23][34] = 8'hb2;
frames[9][23][35] = 8'h6d;
frames[9][23][36] = 8'hb6;
frames[9][23][37] = 8'h92;
frames[9][23][38] = 8'h48;
frames[9][23][39] = 8'hb6;
frames[9][24][0] = 8'hd6;
frames[9][24][1] = 8'hb1;
frames[9][24][2] = 8'had;
frames[9][24][3] = 8'h8c;
frames[9][24][4] = 8'hac;
frames[9][24][5] = 8'hac;
frames[9][24][6] = 8'hac;
frames[9][24][7] = 8'h8c;
frames[9][24][8] = 8'h88;
frames[9][24][9] = 8'h88;
frames[9][24][10] = 8'hac;
frames[9][24][11] = 8'hac;
frames[9][24][12] = 8'hac;
frames[9][24][13] = 8'h88;
frames[9][24][14] = 8'h68;
frames[9][24][15] = 8'h64;
frames[9][24][16] = 8'h48;
frames[9][24][17] = 8'h24;
frames[9][24][18] = 8'h24;
frames[9][24][19] = 8'h44;
frames[9][24][20] = 8'h44;
frames[9][24][21] = 8'h44;
frames[9][24][22] = 8'h44;
frames[9][24][23] = 8'h8d;
frames[9][24][24] = 8'hd6;
frames[9][24][25] = 8'hd6;
frames[9][24][26] = 8'hd6;
frames[9][24][27] = 8'hd6;
frames[9][24][28] = 8'hd6;
frames[9][24][29] = 8'hd6;
frames[9][24][30] = 8'hda;
frames[9][24][31] = 8'hda;
frames[9][24][32] = 8'hb6;
frames[9][24][33] = 8'h8d;
frames[9][24][34] = 8'h24;
frames[9][24][35] = 8'h49;
frames[9][24][36] = 8'hb6;
frames[9][24][37] = 8'h92;
frames[9][24][38] = 8'h49;
frames[9][24][39] = 8'h6d;
frames[9][25][0] = 8'hb1;
frames[9][25][1] = 8'hb1;
frames[9][25][2] = 8'hac;
frames[9][25][3] = 8'hac;
frames[9][25][4] = 8'hac;
frames[9][25][5] = 8'hac;
frames[9][25][6] = 8'hac;
frames[9][25][7] = 8'hac;
frames[9][25][8] = 8'hac;
frames[9][25][9] = 8'hac;
frames[9][25][10] = 8'hb0;
frames[9][25][11] = 8'hac;
frames[9][25][12] = 8'hac;
frames[9][25][13] = 8'h88;
frames[9][25][14] = 8'h68;
frames[9][25][15] = 8'h64;
frames[9][25][16] = 8'h44;
frames[9][25][17] = 8'h44;
frames[9][25][18] = 8'h24;
frames[9][25][19] = 8'h44;
frames[9][25][20] = 8'h24;
frames[9][25][21] = 8'h24;
frames[9][25][22] = 8'h24;
frames[9][25][23] = 8'h24;
frames[9][25][24] = 8'h44;
frames[9][25][25] = 8'h6d;
frames[9][25][26] = 8'h8d;
frames[9][25][27] = 8'h91;
frames[9][25][28] = 8'h91;
frames[9][25][29] = 8'h91;
frames[9][25][30] = 8'h8d;
frames[9][25][31] = 8'h69;
frames[9][25][32] = 8'h24;
frames[9][25][33] = 8'h24;
frames[9][25][34] = 8'h44;
frames[9][25][35] = 8'h91;
frames[9][25][36] = 8'hb6;
frames[9][25][37] = 8'h96;
frames[9][25][38] = 8'h49;
frames[9][25][39] = 8'h6d;
frames[9][26][0] = 8'hb1;
frames[9][26][1] = 8'hb1;
frames[9][26][2] = 8'hac;
frames[9][26][3] = 8'hac;
frames[9][26][4] = 8'hac;
frames[9][26][5] = 8'hac;
frames[9][26][6] = 8'hac;
frames[9][26][7] = 8'hac;
frames[9][26][8] = 8'hb0;
frames[9][26][9] = 8'hb0;
frames[9][26][10] = 8'hb0;
frames[9][26][11] = 8'hac;
frames[9][26][12] = 8'hac;
frames[9][26][13] = 8'h88;
frames[9][26][14] = 8'h68;
frames[9][26][15] = 8'h64;
frames[9][26][16] = 8'h44;
frames[9][26][17] = 8'h44;
frames[9][26][18] = 8'h48;
frames[9][26][19] = 8'h48;
frames[9][26][20] = 8'h48;
frames[9][26][21] = 8'h48;
frames[9][26][22] = 8'h48;
frames[9][26][23] = 8'h48;
frames[9][26][24] = 8'h44;
frames[9][26][25] = 8'h44;
frames[9][26][26] = 8'h48;
frames[9][26][27] = 8'h69;
frames[9][26][28] = 8'h69;
frames[9][26][29] = 8'h6d;
frames[9][26][30] = 8'h6d;
frames[9][26][31] = 8'h6d;
frames[9][26][32] = 8'h8d;
frames[9][26][33] = 8'h91;
frames[9][26][34] = 8'h92;
frames[9][26][35] = 8'h92;
frames[9][26][36] = 8'h6d;
frames[9][26][37] = 8'h49;
frames[9][26][38] = 8'h48;
frames[9][26][39] = 8'h91;
frames[9][27][0] = 8'hb1;
frames[9][27][1] = 8'hb1;
frames[9][27][2] = 8'hb1;
frames[9][27][3] = 8'hb1;
frames[9][27][4] = 8'hac;
frames[9][27][5] = 8'hac;
frames[9][27][6] = 8'hac;
frames[9][27][7] = 8'hb0;
frames[9][27][8] = 8'hb0;
frames[9][27][9] = 8'hb0;
frames[9][27][10] = 8'hac;
frames[9][27][11] = 8'hac;
frames[9][27][12] = 8'h8c;
frames[9][27][13] = 8'h88;
frames[9][27][14] = 8'h68;
frames[9][27][15] = 8'h64;
frames[9][27][16] = 8'h44;
frames[9][27][17] = 8'h44;
frames[9][27][18] = 8'h44;
frames[9][27][19] = 8'h44;
frames[9][27][20] = 8'h44;
frames[9][27][21] = 8'h44;
frames[9][27][22] = 8'h44;
frames[9][27][23] = 8'h44;
frames[9][27][24] = 8'h44;
frames[9][27][25] = 8'h44;
frames[9][27][26] = 8'h44;
frames[9][27][27] = 8'h44;
frames[9][27][28] = 8'h44;
frames[9][27][29] = 8'h44;
frames[9][27][30] = 8'h44;
frames[9][27][31] = 8'h44;
frames[9][27][32] = 8'h44;
frames[9][27][33] = 8'h44;
frames[9][27][34] = 8'h44;
frames[9][27][35] = 8'h44;
frames[9][27][36] = 8'h44;
frames[9][27][37] = 8'h44;
frames[9][27][38] = 8'h68;
frames[9][27][39] = 8'hb1;
frames[9][28][0] = 8'hb1;
frames[9][28][1] = 8'hb1;
frames[9][28][2] = 8'hd1;
frames[9][28][3] = 8'hb1;
frames[9][28][4] = 8'hb1;
frames[9][28][5] = 8'hb1;
frames[9][28][6] = 8'hac;
frames[9][28][7] = 8'hac;
frames[9][28][8] = 8'hac;
frames[9][28][9] = 8'hac;
frames[9][28][10] = 8'hac;
frames[9][28][11] = 8'hac;
frames[9][28][12] = 8'h8c;
frames[9][28][13] = 8'h88;
frames[9][28][14] = 8'h64;
frames[9][28][15] = 8'h64;
frames[9][28][16] = 8'h64;
frames[9][28][17] = 8'h64;
frames[9][28][18] = 8'h64;
frames[9][28][19] = 8'h64;
frames[9][28][20] = 8'h44;
frames[9][28][21] = 8'h44;
frames[9][28][22] = 8'h44;
frames[9][28][23] = 8'h44;
frames[9][28][24] = 8'h64;
frames[9][28][25] = 8'h44;
frames[9][28][26] = 8'h44;
frames[9][28][27] = 8'h44;
frames[9][28][28] = 8'h44;
frames[9][28][29] = 8'h44;
frames[9][28][30] = 8'h44;
frames[9][28][31] = 8'h44;
frames[9][28][32] = 8'h44;
frames[9][28][33] = 8'h44;
frames[9][28][34] = 8'h44;
frames[9][28][35] = 8'h44;
frames[9][28][36] = 8'h64;
frames[9][28][37] = 8'h64;
frames[9][28][38] = 8'h88;
frames[9][28][39] = 8'hb1;
frames[9][29][0] = 8'hd1;
frames[9][29][1] = 8'hb1;
frames[9][29][2] = 8'hb1;
frames[9][29][3] = 8'hd1;
frames[9][29][4] = 8'hd1;
frames[9][29][5] = 8'hb1;
frames[9][29][6] = 8'hb0;
frames[9][29][7] = 8'hb0;
frames[9][29][8] = 8'hb1;
frames[9][29][9] = 8'had;
frames[9][29][10] = 8'had;
frames[9][29][11] = 8'had;
frames[9][29][12] = 8'hac;
frames[9][29][13] = 8'h88;
frames[9][29][14] = 8'h88;
frames[9][29][15] = 8'h88;
frames[9][29][16] = 8'h88;
frames[9][29][17] = 8'h88;
frames[9][29][18] = 8'h68;
frames[9][29][19] = 8'h64;
frames[9][29][20] = 8'h64;
frames[9][29][21] = 8'h64;
frames[9][29][22] = 8'h64;
frames[9][29][23] = 8'h64;
frames[9][29][24] = 8'h68;
frames[9][29][25] = 8'h64;
frames[9][29][26] = 8'h64;
frames[9][29][27] = 8'h68;
frames[9][29][28] = 8'h68;
frames[9][29][29] = 8'h68;
frames[9][29][30] = 8'h68;
frames[9][29][31] = 8'h68;
frames[9][29][32] = 8'h68;
frames[9][29][33] = 8'h88;
frames[9][29][34] = 8'h88;
frames[9][29][35] = 8'h8c;
frames[9][29][36] = 8'had;
frames[9][29][37] = 8'hb1;
frames[9][29][38] = 8'hd1;
frames[9][29][39] = 8'hd6;
frames[10][0][0] = 8'hda;
frames[10][0][1] = 8'hda;
frames[10][0][2] = 8'hd6;
frames[10][0][3] = 8'hb2;
frames[10][0][4] = 8'h00;
frames[10][0][5] = 8'h00;
frames[10][0][6] = 8'h00;
frames[10][0][7] = 8'h00;
frames[10][0][8] = 8'h00;
frames[10][0][9] = 8'h00;
frames[10][0][10] = 8'h8d;
frames[10][0][11] = 8'hd2;
frames[10][0][12] = 8'hd1;
frames[10][0][13] = 8'hd1;
frames[10][0][14] = 8'hd1;
frames[10][0][15] = 8'hd1;
frames[10][0][16] = 8'had;
frames[10][0][17] = 8'had;
frames[10][0][18] = 8'h44;
frames[10][0][19] = 8'h00;
frames[10][0][20] = 8'h00;
frames[10][0][21] = 8'h00;
frames[10][0][22] = 8'h00;
frames[10][0][23] = 8'h00;
frames[10][0][24] = 8'h00;
frames[10][0][25] = 8'h00;
frames[10][0][26] = 8'h44;
frames[10][0][27] = 8'h64;
frames[10][0][28] = 8'had;
frames[10][0][29] = 8'hd1;
frames[10][0][30] = 8'hd6;
frames[10][0][31] = 8'hd6;
frames[10][0][32] = 8'hd6;
frames[10][0][33] = 8'hd6;
frames[10][0][34] = 8'hb2;
frames[10][0][35] = 8'hd6;
frames[10][0][36] = 8'hd6;
frames[10][0][37] = 8'hb6;
frames[10][0][38] = 8'hda;
frames[10][0][39] = 8'hd6;
frames[10][1][0] = 8'hda;
frames[10][1][1] = 8'hda;
frames[10][1][2] = 8'hda;
frames[10][1][3] = 8'h91;
frames[10][1][4] = 8'h00;
frames[10][1][5] = 8'h00;
frames[10][1][6] = 8'h00;
frames[10][1][7] = 8'h00;
frames[10][1][8] = 8'h00;
frames[10][1][9] = 8'h00;
frames[10][1][10] = 8'h20;
frames[10][1][11] = 8'h8d;
frames[10][1][12] = 8'hd1;
frames[10][1][13] = 8'hd1;
frames[10][1][14] = 8'hd1;
frames[10][1][15] = 8'hd1;
frames[10][1][16] = 8'hd1;
frames[10][1][17] = 8'hd1;
frames[10][1][18] = 8'h8d;
frames[10][1][19] = 8'h20;
frames[10][1][20] = 8'h00;
frames[10][1][21] = 8'h00;
frames[10][1][22] = 8'h00;
frames[10][1][23] = 8'h00;
frames[10][1][24] = 8'h00;
frames[10][1][25] = 8'h20;
frames[10][1][26] = 8'h44;
frames[10][1][27] = 8'h64;
frames[10][1][28] = 8'h8d;
frames[10][1][29] = 8'hd1;
frames[10][1][30] = 8'hd6;
frames[10][1][31] = 8'hd6;
frames[10][1][32] = 8'hd6;
frames[10][1][33] = 8'hd6;
frames[10][1][34] = 8'hb2;
frames[10][1][35] = 8'hd6;
frames[10][1][36] = 8'hdb;
frames[10][1][37] = 8'hda;
frames[10][1][38] = 8'hdb;
frames[10][1][39] = 8'hdb;
frames[10][2][0] = 8'hda;
frames[10][2][1] = 8'hd6;
frames[10][2][2] = 8'hd6;
frames[10][2][3] = 8'h6d;
frames[10][2][4] = 8'h00;
frames[10][2][5] = 8'h00;
frames[10][2][6] = 8'h00;
frames[10][2][7] = 8'h00;
frames[10][2][8] = 8'h00;
frames[10][2][9] = 8'h00;
frames[10][2][10] = 8'h00;
frames[10][2][11] = 8'h24;
frames[10][2][12] = 8'hb1;
frames[10][2][13] = 8'hd1;
frames[10][2][14] = 8'hd1;
frames[10][2][15] = 8'hd1;
frames[10][2][16] = 8'hd1;
frames[10][2][17] = 8'had;
frames[10][2][18] = 8'had;
frames[10][2][19] = 8'h8d;
frames[10][2][20] = 8'h00;
frames[10][2][21] = 8'h00;
frames[10][2][22] = 8'h00;
frames[10][2][23] = 8'h00;
frames[10][2][24] = 8'h00;
frames[10][2][25] = 8'h24;
frames[10][2][26] = 8'h44;
frames[10][2][27] = 8'h64;
frames[10][2][28] = 8'h8d;
frames[10][2][29] = 8'hb1;
frames[10][2][30] = 8'hd6;
frames[10][2][31] = 8'hd6;
frames[10][2][32] = 8'hd6;
frames[10][2][33] = 8'hd6;
frames[10][2][34] = 8'hb2;
frames[10][2][35] = 8'hd6;
frames[10][2][36] = 8'hdb;
frames[10][2][37] = 8'h92;
frames[10][2][38] = 8'hb2;
frames[10][2][39] = 8'hdb;
frames[10][3][0] = 8'hda;
frames[10][3][1] = 8'hd6;
frames[10][3][2] = 8'hd6;
frames[10][3][3] = 8'h44;
frames[10][3][4] = 8'h00;
frames[10][3][5] = 8'h00;
frames[10][3][6] = 8'h00;
frames[10][3][7] = 8'h00;
frames[10][3][8] = 8'h00;
frames[10][3][9] = 8'h00;
frames[10][3][10] = 8'h00;
frames[10][3][11] = 8'h00;
frames[10][3][12] = 8'h64;
frames[10][3][13] = 8'hb2;
frames[10][3][14] = 8'hd1;
frames[10][3][15] = 8'hd1;
frames[10][3][16] = 8'hd1;
frames[10][3][17] = 8'hd1;
frames[10][3][18] = 8'had;
frames[10][3][19] = 8'had;
frames[10][3][20] = 8'h69;
frames[10][3][21] = 8'h20;
frames[10][3][22] = 8'h00;
frames[10][3][23] = 8'h00;
frames[10][3][24] = 8'h20;
frames[10][3][25] = 8'h48;
frames[10][3][26] = 8'h64;
frames[10][3][27] = 8'h64;
frames[10][3][28] = 8'h8d;
frames[10][3][29] = 8'hd1;
frames[10][3][30] = 8'hd6;
frames[10][3][31] = 8'hd6;
frames[10][3][32] = 8'hd6;
frames[10][3][33] = 8'hd6;
frames[10][3][34] = 8'hb2;
frames[10][3][35] = 8'hd6;
frames[10][3][36] = 8'hda;
frames[10][3][37] = 8'hb2;
frames[10][3][38] = 8'hda;
frames[10][3][39] = 8'hfb;
frames[10][4][0] = 8'hda;
frames[10][4][1] = 8'hd6;
frames[10][4][2] = 8'hb6;
frames[10][4][3] = 8'h24;
frames[10][4][4] = 8'h00;
frames[10][4][5] = 8'h00;
frames[10][4][6] = 8'h00;
frames[10][4][7] = 8'h00;
frames[10][4][8] = 8'h00;
frames[10][4][9] = 8'h00;
frames[10][4][10] = 8'h00;
frames[10][4][11] = 8'h00;
frames[10][4][12] = 8'h00;
frames[10][4][13] = 8'h6d;
frames[10][4][14] = 8'hd1;
frames[10][4][15] = 8'hd1;
frames[10][4][16] = 8'hd1;
frames[10][4][17] = 8'hd1;
frames[10][4][18] = 8'hd1;
frames[10][4][19] = 8'had;
frames[10][4][20] = 8'had;
frames[10][4][21] = 8'h89;
frames[10][4][22] = 8'h00;
frames[10][4][23] = 8'h00;
frames[10][4][24] = 8'h20;
frames[10][4][25] = 8'h69;
frames[10][4][26] = 8'h64;
frames[10][4][27] = 8'h64;
frames[10][4][28] = 8'h89;
frames[10][4][29] = 8'had;
frames[10][4][30] = 8'hd6;
frames[10][4][31] = 8'hd6;
frames[10][4][32] = 8'hd6;
frames[10][4][33] = 8'hd6;
frames[10][4][34] = 8'hb2;
frames[10][4][35] = 8'hd6;
frames[10][4][36] = 8'hdb;
frames[10][4][37] = 8'hb6;
frames[10][4][38] = 8'hda;
frames[10][4][39] = 8'hfb;
frames[10][5][0] = 8'hda;
frames[10][5][1] = 8'hda;
frames[10][5][2] = 8'hb6;
frames[10][5][3] = 8'h00;
frames[10][5][4] = 8'h00;
frames[10][5][5] = 8'h00;
frames[10][5][6] = 8'h00;
frames[10][5][7] = 8'h00;
frames[10][5][8] = 8'h00;
frames[10][5][9] = 8'h00;
frames[10][5][10] = 8'h00;
frames[10][5][11] = 8'h00;
frames[10][5][12] = 8'h00;
frames[10][5][13] = 8'h00;
frames[10][5][14] = 8'h8d;
frames[10][5][15] = 8'hd1;
frames[10][5][16] = 8'hd1;
frames[10][5][17] = 8'hd1;
frames[10][5][18] = 8'hd1;
frames[10][5][19] = 8'hd1;
frames[10][5][20] = 8'had;
frames[10][5][21] = 8'hcd;
frames[10][5][22] = 8'h6d;
frames[10][5][23] = 8'h20;
frames[10][5][24] = 8'h20;
frames[10][5][25] = 8'h69;
frames[10][5][26] = 8'h40;
frames[10][5][27] = 8'h69;
frames[10][5][28] = 8'h88;
frames[10][5][29] = 8'h89;
frames[10][5][30] = 8'hd6;
frames[10][5][31] = 8'hd6;
frames[10][5][32] = 8'hd6;
frames[10][5][33] = 8'hd6;
frames[10][5][34] = 8'hb2;
frames[10][5][35] = 8'hd6;
frames[10][5][36] = 8'hd6;
frames[10][5][37] = 8'hda;
frames[10][5][38] = 8'hdb;
frames[10][5][39] = 8'hda;
frames[10][6][0] = 8'hb6;
frames[10][6][1] = 8'hb6;
frames[10][6][2] = 8'h92;
frames[10][6][3] = 8'h28;
frames[10][6][4] = 8'h24;
frames[10][6][5] = 8'h00;
frames[10][6][6] = 8'h00;
frames[10][6][7] = 8'h00;
frames[10][6][8] = 8'h00;
frames[10][6][9] = 8'h00;
frames[10][6][10] = 8'h00;
frames[10][6][11] = 8'h00;
frames[10][6][12] = 8'h00;
frames[10][6][13] = 8'h00;
frames[10][6][14] = 8'h20;
frames[10][6][15] = 8'h6d;
frames[10][6][16] = 8'hd1;
frames[10][6][17] = 8'hd1;
frames[10][6][18] = 8'hd1;
frames[10][6][19] = 8'hd1;
frames[10][6][20] = 8'hd1;
frames[10][6][21] = 8'had;
frames[10][6][22] = 8'hb1;
frames[10][6][23] = 8'h88;
frames[10][6][24] = 8'h44;
frames[10][6][25] = 8'h68;
frames[10][6][26] = 8'h64;
frames[10][6][27] = 8'h89;
frames[10][6][28] = 8'h68;
frames[10][6][29] = 8'hd1;
frames[10][6][30] = 8'hd6;
frames[10][6][31] = 8'hd6;
frames[10][6][32] = 8'hd6;
frames[10][6][33] = 8'hb6;
frames[10][6][34] = 8'hb2;
frames[10][6][35] = 8'hd6;
frames[10][6][36] = 8'hb6;
frames[10][6][37] = 8'h91;
frames[10][6][38] = 8'hd6;
frames[10][6][39] = 8'hd6;
frames[10][7][0] = 8'h71;
frames[10][7][1] = 8'h71;
frames[10][7][2] = 8'h71;
frames[10][7][3] = 8'h72;
frames[10][7][4] = 8'h92;
frames[10][7][5] = 8'h92;
frames[10][7][6] = 8'h6d;
frames[10][7][7] = 8'h24;
frames[10][7][8] = 8'h00;
frames[10][7][9] = 8'h00;
frames[10][7][10] = 8'h00;
frames[10][7][11] = 8'h00;
frames[10][7][12] = 8'h00;
frames[10][7][13] = 8'h00;
frames[10][7][14] = 8'h00;
frames[10][7][15] = 8'h00;
frames[10][7][16] = 8'h68;
frames[10][7][17] = 8'hb1;
frames[10][7][18] = 8'hd1;
frames[10][7][19] = 8'hd1;
frames[10][7][20] = 8'hd1;
frames[10][7][21] = 8'hcd;
frames[10][7][22] = 8'had;
frames[10][7][23] = 8'had;
frames[10][7][24] = 8'h8d;
frames[10][7][25] = 8'h64;
frames[10][7][26] = 8'h64;
frames[10][7][27] = 8'h68;
frames[10][7][28] = 8'h68;
frames[10][7][29] = 8'hb1;
frames[10][7][30] = 8'hb6;
frames[10][7][31] = 8'hb6;
frames[10][7][32] = 8'hb6;
frames[10][7][33] = 8'hb6;
frames[10][7][34] = 8'hb6;
frames[10][7][35] = 8'hd6;
frames[10][7][36] = 8'hb6;
frames[10][7][37] = 8'hb1;
frames[10][7][38] = 8'hb6;
frames[10][7][39] = 8'hd6;
frames[10][8][0] = 8'h91;
frames[10][8][1] = 8'h92;
frames[10][8][2] = 8'hb6;
frames[10][8][3] = 8'hb6;
frames[10][8][4] = 8'hd6;
frames[10][8][5] = 8'hd6;
frames[10][8][6] = 8'hda;
frames[10][8][7] = 8'hb6;
frames[10][8][8] = 8'h6d;
frames[10][8][9] = 8'h20;
frames[10][8][10] = 8'h20;
frames[10][8][11] = 8'h20;
frames[10][8][12] = 8'h20;
frames[10][8][13] = 8'h20;
frames[10][8][14] = 8'h20;
frames[10][8][15] = 8'h20;
frames[10][8][16] = 8'h20;
frames[10][8][17] = 8'h69;
frames[10][8][18] = 8'had;
frames[10][8][19] = 8'hd1;
frames[10][8][20] = 8'hd1;
frames[10][8][21] = 8'hd1;
frames[10][8][22] = 8'had;
frames[10][8][23] = 8'had;
frames[10][8][24] = 8'had;
frames[10][8][25] = 8'h89;
frames[10][8][26] = 8'h44;
frames[10][8][27] = 8'h44;
frames[10][8][28] = 8'h48;
frames[10][8][29] = 8'h48;
frames[10][8][30] = 8'h69;
frames[10][8][31] = 8'h69;
frames[10][8][32] = 8'h49;
frames[10][8][33] = 8'h49;
frames[10][8][34] = 8'h49;
frames[10][8][35] = 8'h8d;
frames[10][8][36] = 8'hdb;
frames[10][8][37] = 8'hdb;
frames[10][8][38] = 8'hfb;
frames[10][8][39] = 8'hfb;
frames[10][9][0] = 8'hd6;
frames[10][9][1] = 8'hd6;
frames[10][9][2] = 8'hd6;
frames[10][9][3] = 8'hb6;
frames[10][9][4] = 8'hb6;
frames[10][9][5] = 8'hb6;
frames[10][9][6] = 8'hb6;
frames[10][9][7] = 8'hd6;
frames[10][9][8] = 8'hb2;
frames[10][9][9] = 8'h6d;
frames[10][9][10] = 8'h44;
frames[10][9][11] = 8'h44;
frames[10][9][12] = 8'h44;
frames[10][9][13] = 8'h44;
frames[10][9][14] = 8'h44;
frames[10][9][15] = 8'h44;
frames[10][9][16] = 8'h44;
frames[10][9][17] = 8'h44;
frames[10][9][18] = 8'h68;
frames[10][9][19] = 8'hb1;
frames[10][9][20] = 8'hd1;
frames[10][9][21] = 8'hd1;
frames[10][9][22] = 8'hd1;
frames[10][9][23] = 8'had;
frames[10][9][24] = 8'had;
frames[10][9][25] = 8'had;
frames[10][9][26] = 8'h8d;
frames[10][9][27] = 8'h8d;
frames[10][9][28] = 8'h8d;
frames[10][9][29] = 8'h6d;
frames[10][9][30] = 8'h44;
frames[10][9][31] = 8'h24;
frames[10][9][32] = 8'h24;
frames[10][9][33] = 8'h20;
frames[10][9][34] = 8'h00;
frames[10][9][35] = 8'h24;
frames[10][9][36] = 8'hfb;
frames[10][9][37] = 8'hff;
frames[10][9][38] = 8'hff;
frames[10][9][39] = 8'hff;
frames[10][10][0] = 8'hd6;
frames[10][10][1] = 8'hd6;
frames[10][10][2] = 8'hd6;
frames[10][10][3] = 8'hd6;
frames[10][10][4] = 8'hd6;
frames[10][10][5] = 8'hd6;
frames[10][10][6] = 8'hb6;
frames[10][10][7] = 8'hb1;
frames[10][10][8] = 8'h91;
frames[10][10][9] = 8'h6d;
frames[10][10][10] = 8'h68;
frames[10][10][11] = 8'h68;
frames[10][10][12] = 8'h68;
frames[10][10][13] = 8'h68;
frames[10][10][14] = 8'h44;
frames[10][10][15] = 8'h44;
frames[10][10][16] = 8'h24;
frames[10][10][17] = 8'h24;
frames[10][10][18] = 8'h24;
frames[10][10][19] = 8'h44;
frames[10][10][20] = 8'had;
frames[10][10][21] = 8'hb1;
frames[10][10][22] = 8'hd1;
frames[10][10][23] = 8'had;
frames[10][10][24] = 8'had;
frames[10][10][25] = 8'had;
frames[10][10][26] = 8'hb1;
frames[10][10][27] = 8'hd6;
frames[10][10][28] = 8'hda;
frames[10][10][29] = 8'hd6;
frames[10][10][30] = 8'hb6;
frames[10][10][31] = 8'h8d;
frames[10][10][32] = 8'h69;
frames[10][10][33] = 8'h69;
frames[10][10][34] = 8'h49;
frames[10][10][35] = 8'h24;
frames[10][10][36] = 8'hd6;
frames[10][10][37] = 8'hff;
frames[10][10][38] = 8'hff;
frames[10][10][39] = 8'hff;
frames[10][11][0] = 8'hd6;
frames[10][11][1] = 8'hd6;
frames[10][11][2] = 8'hd6;
frames[10][11][3] = 8'hd6;
frames[10][11][4] = 8'hd6;
frames[10][11][5] = 8'hd6;
frames[10][11][6] = 8'hb6;
frames[10][11][7] = 8'hb1;
frames[10][11][8] = 8'h8d;
frames[10][11][9] = 8'h6d;
frames[10][11][10] = 8'h68;
frames[10][11][11] = 8'h68;
frames[10][11][12] = 8'h88;
frames[10][11][13] = 8'h68;
frames[10][11][14] = 8'h44;
frames[10][11][15] = 8'h40;
frames[10][11][16] = 8'h24;
frames[10][11][17] = 8'h24;
frames[10][11][18] = 8'h24;
frames[10][11][19] = 8'h24;
frames[10][11][20] = 8'h69;
frames[10][11][21] = 8'hb6;
frames[10][11][22] = 8'hb1;
frames[10][11][23] = 8'hb1;
frames[10][11][24] = 8'had;
frames[10][11][25] = 8'had;
frames[10][11][26] = 8'had;
frames[10][11][27] = 8'hb1;
frames[10][11][28] = 8'hd6;
frames[10][11][29] = 8'hfa;
frames[10][11][30] = 8'hda;
frames[10][11][31] = 8'hd6;
frames[10][11][32] = 8'hb2;
frames[10][11][33] = 8'hb2;
frames[10][11][34] = 8'hb2;
frames[10][11][35] = 8'h49;
frames[10][11][36] = 8'h92;
frames[10][11][37] = 8'hff;
frames[10][11][38] = 8'hff;
frames[10][11][39] = 8'hff;
frames[10][12][0] = 8'hd6;
frames[10][12][1] = 8'hd6;
frames[10][12][2] = 8'hd6;
frames[10][12][3] = 8'hd6;
frames[10][12][4] = 8'hb6;
frames[10][12][5] = 8'hb6;
frames[10][12][6] = 8'hb6;
frames[10][12][7] = 8'hb1;
frames[10][12][8] = 8'h8d;
frames[10][12][9] = 8'h6d;
frames[10][12][10] = 8'h68;
frames[10][12][11] = 8'h88;
frames[10][12][12] = 8'h88;
frames[10][12][13] = 8'h88;
frames[10][12][14] = 8'h44;
frames[10][12][15] = 8'h40;
frames[10][12][16] = 8'h24;
frames[10][12][17] = 8'h24;
frames[10][12][18] = 8'h24;
frames[10][12][19] = 8'h24;
frames[10][12][20] = 8'hb2;
frames[10][12][21] = 8'hda;
frames[10][12][22] = 8'hd1;
frames[10][12][23] = 8'hb1;
frames[10][12][24] = 8'hd1;
frames[10][12][25] = 8'had;
frames[10][12][26] = 8'had;
frames[10][12][27] = 8'had;
frames[10][12][28] = 8'had;
frames[10][12][29] = 8'hd6;
frames[10][12][30] = 8'hfa;
frames[10][12][31] = 8'hd6;
frames[10][12][32] = 8'hd6;
frames[10][12][33] = 8'hd6;
frames[10][12][34] = 8'hb6;
frames[10][12][35] = 8'h6d;
frames[10][12][36] = 8'h6d;
frames[10][12][37] = 8'hff;
frames[10][12][38] = 8'hff;
frames[10][12][39] = 8'hff;
frames[10][13][0] = 8'hd6;
frames[10][13][1] = 8'hd6;
frames[10][13][2] = 8'hb6;
frames[10][13][3] = 8'hb6;
frames[10][13][4] = 8'hb1;
frames[10][13][5] = 8'h91;
frames[10][13][6] = 8'hb2;
frames[10][13][7] = 8'hb1;
frames[10][13][8] = 8'h8d;
frames[10][13][9] = 8'h68;
frames[10][13][10] = 8'h88;
frames[10][13][11] = 8'h8c;
frames[10][13][12] = 8'h88;
frames[10][13][13] = 8'h88;
frames[10][13][14] = 8'h44;
frames[10][13][15] = 8'h40;
frames[10][13][16] = 8'h24;
frames[10][13][17] = 8'h24;
frames[10][13][18] = 8'h24;
frames[10][13][19] = 8'h20;
frames[10][13][20] = 8'h8d;
frames[10][13][21] = 8'hd6;
frames[10][13][22] = 8'hd6;
frames[10][13][23] = 8'hb1;
frames[10][13][24] = 8'hd1;
frames[10][13][25] = 8'hd1;
frames[10][13][26] = 8'hd1;
frames[10][13][27] = 8'had;
frames[10][13][28] = 8'had;
frames[10][13][29] = 8'had;
frames[10][13][30] = 8'hd5;
frames[10][13][31] = 8'hf6;
frames[10][13][32] = 8'hd6;
frames[10][13][33] = 8'hd6;
frames[10][13][34] = 8'hb6;
frames[10][13][35] = 8'h91;
frames[10][13][36] = 8'h69;
frames[10][13][37] = 8'hff;
frames[10][13][38] = 8'hff;
frames[10][13][39] = 8'hff;
frames[10][14][0] = 8'hb6;
frames[10][14][1] = 8'hb2;
frames[10][14][2] = 8'h91;
frames[10][14][3] = 8'h91;
frames[10][14][4] = 8'h8d;
frames[10][14][5] = 8'h6d;
frames[10][14][6] = 8'hb2;
frames[10][14][7] = 8'hb2;
frames[10][14][8] = 8'h68;
frames[10][14][9] = 8'h68;
frames[10][14][10] = 8'h8c;
frames[10][14][11] = 8'h8c;
frames[10][14][12] = 8'h88;
frames[10][14][13] = 8'h88;
frames[10][14][14] = 8'h44;
frames[10][14][15] = 8'h40;
frames[10][14][16] = 8'h24;
frames[10][14][17] = 8'h24;
frames[10][14][18] = 8'h24;
frames[10][14][19] = 8'h20;
frames[10][14][20] = 8'h24;
frames[10][14][21] = 8'h91;
frames[10][14][22] = 8'hd6;
frames[10][14][23] = 8'hb1;
frames[10][14][24] = 8'hd1;
frames[10][14][25] = 8'hd1;
frames[10][14][26] = 8'hd1;
frames[10][14][27] = 8'had;
frames[10][14][28] = 8'had;
frames[10][14][29] = 8'had;
frames[10][14][30] = 8'hb1;
frames[10][14][31] = 8'hf6;
frames[10][14][32] = 8'hda;
frames[10][14][33] = 8'hd6;
frames[10][14][34] = 8'hb6;
frames[10][14][35] = 8'h92;
frames[10][14][36] = 8'h49;
frames[10][14][37] = 8'hdb;
frames[10][14][38] = 8'hff;
frames[10][14][39] = 8'hff;
frames[10][15][0] = 8'h91;
frames[10][15][1] = 8'hb2;
frames[10][15][2] = 8'hb2;
frames[10][15][3] = 8'hb6;
frames[10][15][4] = 8'hb2;
frames[10][15][5] = 8'h8d;
frames[10][15][6] = 8'h91;
frames[10][15][7] = 8'hb1;
frames[10][15][8] = 8'h68;
frames[10][15][9] = 8'h68;
frames[10][15][10] = 8'h8c;
frames[10][15][11] = 8'h8d;
frames[10][15][12] = 8'h8c;
frames[10][15][13] = 8'h68;
frames[10][15][14] = 8'h44;
frames[10][15][15] = 8'h40;
frames[10][15][16] = 8'h24;
frames[10][15][17] = 8'h24;
frames[10][15][18] = 8'h24;
frames[10][15][19] = 8'h24;
frames[10][15][20] = 8'h24;
frames[10][15][21] = 8'h24;
frames[10][15][22] = 8'h8d;
frames[10][15][23] = 8'hb1;
frames[10][15][24] = 8'hd1;
frames[10][15][25] = 8'hd1;
frames[10][15][26] = 8'hd1;
frames[10][15][27] = 8'hd1;
frames[10][15][28] = 8'had;
frames[10][15][29] = 8'had;
frames[10][15][30] = 8'had;
frames[10][15][31] = 8'hd6;
frames[10][15][32] = 8'hb6;
frames[10][15][33] = 8'h6d;
frames[10][15][34] = 8'h92;
frames[10][15][35] = 8'hb6;
frames[10][15][36] = 8'h49;
frames[10][15][37] = 8'hb6;
frames[10][15][38] = 8'hff;
frames[10][15][39] = 8'hff;
frames[10][16][0] = 8'h91;
frames[10][16][1] = 8'h8d;
frames[10][16][2] = 8'h91;
frames[10][16][3] = 8'hd6;
frames[10][16][4] = 8'hd6;
frames[10][16][5] = 8'hda;
frames[10][16][6] = 8'hd6;
frames[10][16][7] = 8'h8d;
frames[10][16][8] = 8'h68;
frames[10][16][9] = 8'h8d;
frames[10][16][10] = 8'h8d;
frames[10][16][11] = 8'h8d;
frames[10][16][12] = 8'h88;
frames[10][16][13] = 8'h68;
frames[10][16][14] = 8'h44;
frames[10][16][15] = 8'h44;
frames[10][16][16] = 8'h44;
frames[10][16][17] = 8'h24;
frames[10][16][18] = 8'h24;
frames[10][16][19] = 8'h24;
frames[10][16][20] = 8'h24;
frames[10][16][21] = 8'h24;
frames[10][16][22] = 8'h24;
frames[10][16][23] = 8'h44;
frames[10][16][24] = 8'had;
frames[10][16][25] = 8'had;
frames[10][16][26] = 8'hcd;
frames[10][16][27] = 8'hd1;
frames[10][16][28] = 8'hcd;
frames[10][16][29] = 8'h89;
frames[10][16][30] = 8'hb1;
frames[10][16][31] = 8'had;
frames[10][16][32] = 8'h69;
frames[10][16][33] = 8'h91;
frames[10][16][34] = 8'hb6;
frames[10][16][35] = 8'hb6;
frames[10][16][36] = 8'h69;
frames[10][16][37] = 8'h92;
frames[10][16][38] = 8'hff;
frames[10][16][39] = 8'hff;
frames[10][17][0] = 8'h8d;
frames[10][17][1] = 8'hb1;
frames[10][17][2] = 8'hb5;
frames[10][17][3] = 8'hd6;
frames[10][17][4] = 8'hd6;
frames[10][17][5] = 8'hd6;
frames[10][17][6] = 8'hd6;
frames[10][17][7] = 8'hd5;
frames[10][17][8] = 8'hb1;
frames[10][17][9] = 8'h8d;
frames[10][17][10] = 8'h8d;
frames[10][17][11] = 8'h8d;
frames[10][17][12] = 8'h88;
frames[10][17][13] = 8'h68;
frames[10][17][14] = 8'h44;
frames[10][17][15] = 8'h44;
frames[10][17][16] = 8'h44;
frames[10][17][17] = 8'h24;
frames[10][17][18] = 8'h24;
frames[10][17][19] = 8'h24;
frames[10][17][20] = 8'h24;
frames[10][17][21] = 8'h44;
frames[10][17][22] = 8'h44;
frames[10][17][23] = 8'h44;
frames[10][17][24] = 8'h64;
frames[10][17][25] = 8'h8d;
frames[10][17][26] = 8'hcd;
frames[10][17][27] = 8'had;
frames[10][17][28] = 8'hd1;
frames[10][17][29] = 8'had;
frames[10][17][30] = 8'had;
frames[10][17][31] = 8'had;
frames[10][17][32] = 8'h92;
frames[10][17][33] = 8'hb2;
frames[10][17][34] = 8'hb6;
frames[10][17][35] = 8'hb6;
frames[10][17][36] = 8'h6d;
frames[10][17][37] = 8'h6d;
frames[10][17][38] = 8'hff;
frames[10][17][39] = 8'hff;
frames[10][18][0] = 8'hb1;
frames[10][18][1] = 8'hd6;
frames[10][18][2] = 8'hd5;
frames[10][18][3] = 8'hd6;
frames[10][18][4] = 8'hd5;
frames[10][18][5] = 8'hd5;
frames[10][18][6] = 8'hd5;
frames[10][18][7] = 8'hd5;
frames[10][18][8] = 8'hd5;
frames[10][18][9] = 8'hb1;
frames[10][18][10] = 8'hb1;
frames[10][18][11] = 8'h8c;
frames[10][18][12] = 8'h88;
frames[10][18][13] = 8'h68;
frames[10][18][14] = 8'h44;
frames[10][18][15] = 8'h44;
frames[10][18][16] = 8'h44;
frames[10][18][17] = 8'h24;
frames[10][18][18] = 8'h24;
frames[10][18][19] = 8'h24;
frames[10][18][20] = 8'h44;
frames[10][18][21] = 8'h44;
frames[10][18][22] = 8'h44;
frames[10][18][23] = 8'h49;
frames[10][18][24] = 8'h8d;
frames[10][18][25] = 8'hb1;
frames[10][18][26] = 8'had;
frames[10][18][27] = 8'had;
frames[10][18][28] = 8'had;
frames[10][18][29] = 8'hd1;
frames[10][18][30] = 8'had;
frames[10][18][31] = 8'had;
frames[10][18][32] = 8'h8d;
frames[10][18][33] = 8'hb2;
frames[10][18][34] = 8'hb6;
frames[10][18][35] = 8'hb6;
frames[10][18][36] = 8'h8d;
frames[10][18][37] = 8'h69;
frames[10][18][38] = 8'hfb;
frames[10][18][39] = 8'hff;
frames[10][19][0] = 8'h8d;
frames[10][19][1] = 8'hd5;
frames[10][19][2] = 8'hda;
frames[10][19][3] = 8'hd6;
frames[10][19][4] = 8'hda;
frames[10][19][5] = 8'hd6;
frames[10][19][6] = 8'hd5;
frames[10][19][7] = 8'hd5;
frames[10][19][8] = 8'hd5;
frames[10][19][9] = 8'hb1;
frames[10][19][10] = 8'hb1;
frames[10][19][11] = 8'h8c;
frames[10][19][12] = 8'h88;
frames[10][19][13] = 8'h68;
frames[10][19][14] = 8'h44;
frames[10][19][15] = 8'h44;
frames[10][19][16] = 8'h44;
frames[10][19][17] = 8'h24;
frames[10][19][18] = 8'h24;
frames[10][19][19] = 8'h24;
frames[10][19][20] = 8'h44;
frames[10][19][21] = 8'h44;
frames[10][19][22] = 8'h8d;
frames[10][19][23] = 8'hd6;
frames[10][19][24] = 8'hd6;
frames[10][19][25] = 8'hd6;
frames[10][19][26] = 8'hb1;
frames[10][19][27] = 8'had;
frames[10][19][28] = 8'had;
frames[10][19][29] = 8'hcd;
frames[10][19][30] = 8'had;
frames[10][19][31] = 8'had;
frames[10][19][32] = 8'hb1;
frames[10][19][33] = 8'hb1;
frames[10][19][34] = 8'hb2;
frames[10][19][35] = 8'hb6;
frames[10][19][36] = 8'h92;
frames[10][19][37] = 8'h49;
frames[10][19][38] = 8'hda;
frames[10][19][39] = 8'hff;
frames[10][20][0] = 8'hb1;
frames[10][20][1] = 8'hb1;
frames[10][20][2] = 8'hd5;
frames[10][20][3] = 8'hd5;
frames[10][20][4] = 8'hd5;
frames[10][20][5] = 8'hd5;
frames[10][20][6] = 8'hd5;
frames[10][20][7] = 8'hb5;
frames[10][20][8] = 8'hb5;
frames[10][20][9] = 8'hd5;
frames[10][20][10] = 8'hd1;
frames[10][20][11] = 8'h8c;
frames[10][20][12] = 8'h88;
frames[10][20][13] = 8'h88;
frames[10][20][14] = 8'h64;
frames[10][20][15] = 8'h44;
frames[10][20][16] = 8'h48;
frames[10][20][17] = 8'h24;
frames[10][20][18] = 8'h24;
frames[10][20][19] = 8'h24;
frames[10][20][20] = 8'h44;
frames[10][20][21] = 8'h69;
frames[10][20][22] = 8'hd6;
frames[10][20][23] = 8'hd6;
frames[10][20][24] = 8'hd6;
frames[10][20][25] = 8'hd6;
frames[10][20][26] = 8'hd2;
frames[10][20][27] = 8'had;
frames[10][20][28] = 8'had;
frames[10][20][29] = 8'had;
frames[10][20][30] = 8'had;
frames[10][20][31] = 8'had;
frames[10][20][32] = 8'hb1;
frames[10][20][33] = 8'hd6;
frames[10][20][34] = 8'hb6;
frames[10][20][35] = 8'hb6;
frames[10][20][36] = 8'h92;
frames[10][20][37] = 8'h49;
frames[10][20][38] = 8'hb6;
frames[10][20][39] = 8'hff;
frames[10][21][0] = 8'hb1;
frames[10][21][1] = 8'hb1;
frames[10][21][2] = 8'hd6;
frames[10][21][3] = 8'hd6;
frames[10][21][4] = 8'hd6;
frames[10][21][5] = 8'hd6;
frames[10][21][6] = 8'hd5;
frames[10][21][7] = 8'hd5;
frames[10][21][8] = 8'hd5;
frames[10][21][9] = 8'hd5;
frames[10][21][10] = 8'had;
frames[10][21][11] = 8'h8c;
frames[10][21][12] = 8'h8c;
frames[10][21][13] = 8'h88;
frames[10][21][14] = 8'h64;
frames[10][21][15] = 8'h44;
frames[10][21][16] = 8'h48;
frames[10][21][17] = 8'h24;
frames[10][21][18] = 8'h24;
frames[10][21][19] = 8'h24;
frames[10][21][20] = 8'h24;
frames[10][21][21] = 8'h91;
frames[10][21][22] = 8'hd6;
frames[10][21][23] = 8'hb6;
frames[10][21][24] = 8'hb6;
frames[10][21][25] = 8'hb6;
frames[10][21][26] = 8'hd6;
frames[10][21][27] = 8'hb1;
frames[10][21][28] = 8'had;
frames[10][21][29] = 8'hd1;
frames[10][21][30] = 8'had;
frames[10][21][31] = 8'had;
frames[10][21][32] = 8'hb1;
frames[10][21][33] = 8'hd5;
frames[10][21][34] = 8'hd6;
frames[10][21][35] = 8'hd6;
frames[10][21][36] = 8'hb6;
frames[10][21][37] = 8'h49;
frames[10][21][38] = 8'h91;
frames[10][21][39] = 8'hff;
frames[10][22][0] = 8'hd6;
frames[10][22][1] = 8'hb1;
frames[10][22][2] = 8'hb1;
frames[10][22][3] = 8'hd5;
frames[10][22][4] = 8'hd6;
frames[10][22][5] = 8'hd6;
frames[10][22][6] = 8'hd5;
frames[10][22][7] = 8'hd5;
frames[10][22][8] = 8'hd1;
frames[10][22][9] = 8'hb1;
frames[10][22][10] = 8'hac;
frames[10][22][11] = 8'hac;
frames[10][22][12] = 8'hac;
frames[10][22][13] = 8'h88;
frames[10][22][14] = 8'h64;
frames[10][22][15] = 8'h44;
frames[10][22][16] = 8'h48;
frames[10][22][17] = 8'h24;
frames[10][22][18] = 8'h24;
frames[10][22][19] = 8'h24;
frames[10][22][20] = 8'h24;
frames[10][22][21] = 8'h8d;
frames[10][22][22] = 8'hd6;
frames[10][22][23] = 8'hb6;
frames[10][22][24] = 8'hb6;
frames[10][22][25] = 8'hb6;
frames[10][22][26] = 8'hb5;
frames[10][22][27] = 8'hd6;
frames[10][22][28] = 8'hb1;
frames[10][22][29] = 8'hb1;
frames[10][22][30] = 8'had;
frames[10][22][31] = 8'hd5;
frames[10][22][32] = 8'hd5;
frames[10][22][33] = 8'hd6;
frames[10][22][34] = 8'hd6;
frames[10][22][35] = 8'hb6;
frames[10][22][36] = 8'hb6;
frames[10][22][37] = 8'h6d;
frames[10][22][38] = 8'h6d;
frames[10][22][39] = 8'hff;
frames[10][23][0] = 8'hd6;
frames[10][23][1] = 8'hb1;
frames[10][23][2] = 8'h8c;
frames[10][23][3] = 8'hb1;
frames[10][23][4] = 8'hd1;
frames[10][23][5] = 8'hd5;
frames[10][23][6] = 8'hd1;
frames[10][23][7] = 8'hb1;
frames[10][23][8] = 8'hac;
frames[10][23][9] = 8'hac;
frames[10][23][10] = 8'hac;
frames[10][23][11] = 8'hac;
frames[10][23][12] = 8'h88;
frames[10][23][13] = 8'h88;
frames[10][23][14] = 8'h64;
frames[10][23][15] = 8'h44;
frames[10][23][16] = 8'h48;
frames[10][23][17] = 8'h24;
frames[10][23][18] = 8'h24;
frames[10][23][19] = 8'h24;
frames[10][23][20] = 8'h24;
frames[10][23][21] = 8'h49;
frames[10][23][22] = 8'hb6;
frames[10][23][23] = 8'hb6;
frames[10][23][24] = 8'hb6;
frames[10][23][25] = 8'hb2;
frames[10][23][26] = 8'hb1;
frames[10][23][27] = 8'hd6;
frames[10][23][28] = 8'hd5;
frames[10][23][29] = 8'hd5;
frames[10][23][30] = 8'hd5;
frames[10][23][31] = 8'hfa;
frames[10][23][32] = 8'hd6;
frames[10][23][33] = 8'hd6;
frames[10][23][34] = 8'h6d;
frames[10][23][35] = 8'h8d;
frames[10][23][36] = 8'hb6;
frames[10][23][37] = 8'h6d;
frames[10][23][38] = 8'h49;
frames[10][23][39] = 8'hdb;
frames[10][24][0] = 8'hd1;
frames[10][24][1] = 8'had;
frames[10][24][2] = 8'hac;
frames[10][24][3] = 8'hac;
frames[10][24][4] = 8'hac;
frames[10][24][5] = 8'hac;
frames[10][24][6] = 8'h8c;
frames[10][24][7] = 8'h88;
frames[10][24][8] = 8'hac;
frames[10][24][9] = 8'hac;
frames[10][24][10] = 8'hac;
frames[10][24][11] = 8'hac;
frames[10][24][12] = 8'h88;
frames[10][24][13] = 8'h88;
frames[10][24][14] = 8'h64;
frames[10][24][15] = 8'h44;
frames[10][24][16] = 8'h44;
frames[10][24][17] = 8'h24;
frames[10][24][18] = 8'h24;
frames[10][24][19] = 8'h24;
frames[10][24][20] = 8'h24;
frames[10][24][21] = 8'h24;
frames[10][24][22] = 8'h48;
frames[10][24][23] = 8'h8d;
frames[10][24][24] = 8'hb1;
frames[10][24][25] = 8'hb1;
frames[10][24][26] = 8'hb1;
frames[10][24][27] = 8'hb1;
frames[10][24][28] = 8'hb1;
frames[10][24][29] = 8'hb1;
frames[10][24][30] = 8'hb1;
frames[10][24][31] = 8'hd6;
frames[10][24][32] = 8'hb2;
frames[10][24][33] = 8'h48;
frames[10][24][34] = 8'h24;
frames[10][24][35] = 8'h91;
frames[10][24][36] = 8'hb6;
frames[10][24][37] = 8'h92;
frames[10][24][38] = 8'h44;
frames[10][24][39] = 8'hb6;
frames[10][25][0] = 8'hb1;
frames[10][25][1] = 8'had;
frames[10][25][2] = 8'hac;
frames[10][25][3] = 8'hac;
frames[10][25][4] = 8'hac;
frames[10][25][5] = 8'hac;
frames[10][25][6] = 8'hac;
frames[10][25][7] = 8'hac;
frames[10][25][8] = 8'hac;
frames[10][25][9] = 8'hac;
frames[10][25][10] = 8'hac;
frames[10][25][11] = 8'hac;
frames[10][25][12] = 8'h88;
frames[10][25][13] = 8'h88;
frames[10][25][14] = 8'h64;
frames[10][25][15] = 8'h44;
frames[10][25][16] = 8'h44;
frames[10][25][17] = 8'h24;
frames[10][25][18] = 8'h24;
frames[10][25][19] = 8'h24;
frames[10][25][20] = 8'h24;
frames[10][25][21] = 8'h24;
frames[10][25][22] = 8'h24;
frames[10][25][23] = 8'h24;
frames[10][25][24] = 8'h44;
frames[10][25][25] = 8'h48;
frames[10][25][26] = 8'h68;
frames[10][25][27] = 8'h68;
frames[10][25][28] = 8'h68;
frames[10][25][29] = 8'h69;
frames[10][25][30] = 8'h68;
frames[10][25][31] = 8'h44;
frames[10][25][32] = 8'h48;
frames[10][25][33] = 8'h44;
frames[10][25][34] = 8'h6d;
frames[10][25][35] = 8'hb6;
frames[10][25][36] = 8'hb6;
frames[10][25][37] = 8'h92;
frames[10][25][38] = 8'h49;
frames[10][25][39] = 8'hb2;
frames[10][26][0] = 8'hb1;
frames[10][26][1] = 8'hb1;
frames[10][26][2] = 8'hb1;
frames[10][26][3] = 8'hb1;
frames[10][26][4] = 8'hb1;
frames[10][26][5] = 8'hac;
frames[10][26][6] = 8'hac;
frames[10][26][7] = 8'hac;
frames[10][26][8] = 8'hac;
frames[10][26][9] = 8'hac;
frames[10][26][10] = 8'hac;
frames[10][26][11] = 8'hac;
frames[10][26][12] = 8'h88;
frames[10][26][13] = 8'h68;
frames[10][26][14] = 8'h64;
frames[10][26][15] = 8'h64;
frames[10][26][16] = 8'h44;
frames[10][26][17] = 8'h44;
frames[10][26][18] = 8'h48;
frames[10][26][19] = 8'h48;
frames[10][26][20] = 8'h48;
frames[10][26][21] = 8'h44;
frames[10][26][22] = 8'h44;
frames[10][26][23] = 8'h44;
frames[10][26][24] = 8'h44;
frames[10][26][25] = 8'h44;
frames[10][26][26] = 8'h44;
frames[10][26][27] = 8'h44;
frames[10][26][28] = 8'h44;
frames[10][26][29] = 8'h44;
frames[10][26][30] = 8'h44;
frames[10][26][31] = 8'h48;
frames[10][26][32] = 8'h6d;
frames[10][26][33] = 8'h8d;
frames[10][26][34] = 8'h8d;
frames[10][26][35] = 8'h6d;
frames[10][26][36] = 8'h69;
frames[10][26][37] = 8'h49;
frames[10][26][38] = 8'h69;
frames[10][26][39] = 8'hd6;
frames[10][27][0] = 8'hb1;
frames[10][27][1] = 8'hb1;
frames[10][27][2] = 8'hd1;
frames[10][27][3] = 8'hb1;
frames[10][27][4] = 8'hd1;
frames[10][27][5] = 8'hb1;
frames[10][27][6] = 8'had;
frames[10][27][7] = 8'had;
frames[10][27][8] = 8'had;
frames[10][27][9] = 8'had;
frames[10][27][10] = 8'had;
frames[10][27][11] = 8'h8c;
frames[10][27][12] = 8'h88;
frames[10][27][13] = 8'h68;
frames[10][27][14] = 8'h64;
frames[10][27][15] = 8'h64;
frames[10][27][16] = 8'h44;
frames[10][27][17] = 8'h44;
frames[10][27][18] = 8'h44;
frames[10][27][19] = 8'h44;
frames[10][27][20] = 8'h44;
frames[10][27][21] = 8'h44;
frames[10][27][22] = 8'h44;
frames[10][27][23] = 8'h44;
frames[10][27][24] = 8'h44;
frames[10][27][25] = 8'h44;
frames[10][27][26] = 8'h44;
frames[10][27][27] = 8'h44;
frames[10][27][28] = 8'h44;
frames[10][27][29] = 8'h44;
frames[10][27][30] = 8'h44;
frames[10][27][31] = 8'h44;
frames[10][27][32] = 8'h44;
frames[10][27][33] = 8'h44;
frames[10][27][34] = 8'h44;
frames[10][27][35] = 8'h44;
frames[10][27][36] = 8'h44;
frames[10][27][37] = 8'h44;
frames[10][27][38] = 8'h8d;
frames[10][27][39] = 8'hd6;
frames[10][28][0] = 8'hb1;
frames[10][28][1] = 8'hb1;
frames[10][28][2] = 8'hb1;
frames[10][28][3] = 8'hd5;
frames[10][28][4] = 8'hd1;
frames[10][28][5] = 8'hb1;
frames[10][28][6] = 8'hb1;
frames[10][28][7] = 8'hb1;
frames[10][28][8] = 8'hb1;
frames[10][28][9] = 8'had;
frames[10][28][10] = 8'had;
frames[10][28][11] = 8'h8c;
frames[10][28][12] = 8'h88;
frames[10][28][13] = 8'h68;
frames[10][28][14] = 8'h64;
frames[10][28][15] = 8'h64;
frames[10][28][16] = 8'h64;
frames[10][28][17] = 8'h64;
frames[10][28][18] = 8'h64;
frames[10][28][19] = 8'h64;
frames[10][28][20] = 8'h44;
frames[10][28][21] = 8'h44;
frames[10][28][22] = 8'h44;
frames[10][28][23] = 8'h64;
frames[10][28][24] = 8'h44;
frames[10][28][25] = 8'h44;
frames[10][28][26] = 8'h44;
frames[10][28][27] = 8'h44;
frames[10][28][28] = 8'h44;
frames[10][28][29] = 8'h44;
frames[10][28][30] = 8'h44;
frames[10][28][31] = 8'h44;
frames[10][28][32] = 8'h44;
frames[10][28][33] = 8'h64;
frames[10][28][34] = 8'h64;
frames[10][28][35] = 8'h64;
frames[10][28][36] = 8'h64;
frames[10][28][37] = 8'h68;
frames[10][28][38] = 8'h8d;
frames[10][28][39] = 8'hd6;
frames[10][29][0] = 8'hb1;
frames[10][29][1] = 8'hb1;
frames[10][29][2] = 8'hb1;
frames[10][29][3] = 8'hd5;
frames[10][29][4] = 8'hd5;
frames[10][29][5] = 8'hb1;
frames[10][29][6] = 8'hb1;
frames[10][29][7] = 8'hb1;
frames[10][29][8] = 8'hb1;
frames[10][29][9] = 8'had;
frames[10][29][10] = 8'hac;
frames[10][29][11] = 8'h8c;
frames[10][29][12] = 8'h88;
frames[10][29][13] = 8'h68;
frames[10][29][14] = 8'h64;
frames[10][29][15] = 8'h68;
frames[10][29][16] = 8'h88;
frames[10][29][17] = 8'h88;
frames[10][29][18] = 8'h68;
frames[10][29][19] = 8'h68;
frames[10][29][20] = 8'h64;
frames[10][29][21] = 8'h64;
frames[10][29][22] = 8'h64;
frames[10][29][23] = 8'h68;
frames[10][29][24] = 8'h68;
frames[10][29][25] = 8'h68;
frames[10][29][26] = 8'h68;
frames[10][29][27] = 8'h68;
frames[10][29][28] = 8'h88;
frames[10][29][29] = 8'h88;
frames[10][29][30] = 8'h88;
frames[10][29][31] = 8'h88;
frames[10][29][32] = 8'h88;
frames[10][29][33] = 8'h8c;
frames[10][29][34] = 8'h8c;
frames[10][29][35] = 8'had;
frames[10][29][36] = 8'hb1;
frames[10][29][37] = 8'hd1;
frames[10][29][38] = 8'hd6;
frames[10][29][39] = 8'hfa;
frames[11][0][0] = 8'h68;
frames[11][0][1] = 8'h64;
frames[11][0][2] = 8'h64;
frames[11][0][3] = 8'h84;
frames[11][0][4] = 8'h84;
frames[11][0][5] = 8'h88;
frames[11][0][6] = 8'h89;
frames[11][0][7] = 8'h89;
frames[11][0][8] = 8'h89;
frames[11][0][9] = 8'h89;
frames[11][0][10] = 8'ha9;
frames[11][0][11] = 8'had;
frames[11][0][12] = 8'had;
frames[11][0][13] = 8'had;
frames[11][0][14] = 8'had;
frames[11][0][15] = 8'had;
frames[11][0][16] = 8'had;
frames[11][0][17] = 8'had;
frames[11][0][18] = 8'had;
frames[11][0][19] = 8'had;
frames[11][0][20] = 8'had;
frames[11][0][21] = 8'h8d;
frames[11][0][22] = 8'had;
frames[11][0][23] = 8'had;
frames[11][0][24] = 8'had;
frames[11][0][25] = 8'h89;
frames[11][0][26] = 8'h40;
frames[11][0][27] = 8'h40;
frames[11][0][28] = 8'h40;
frames[11][0][29] = 8'h64;
frames[11][0][30] = 8'h84;
frames[11][0][31] = 8'h88;
frames[11][0][32] = 8'h8d;
frames[11][0][33] = 8'h44;
frames[11][0][34] = 8'h24;
frames[11][0][35] = 8'h24;
frames[11][0][36] = 8'h24;
frames[11][0][37] = 8'h6d;
frames[11][0][38] = 8'h6d;
frames[11][0][39] = 8'h69;
frames[11][1][0] = 8'h00;
frames[11][1][1] = 8'h20;
frames[11][1][2] = 8'h40;
frames[11][1][3] = 8'h44;
frames[11][1][4] = 8'h64;
frames[11][1][5] = 8'h64;
frames[11][1][6] = 8'h64;
frames[11][1][7] = 8'h68;
frames[11][1][8] = 8'h68;
frames[11][1][9] = 8'h88;
frames[11][1][10] = 8'h88;
frames[11][1][11] = 8'h89;
frames[11][1][12] = 8'had;
frames[11][1][13] = 8'had;
frames[11][1][14] = 8'had;
frames[11][1][15] = 8'had;
frames[11][1][16] = 8'had;
frames[11][1][17] = 8'had;
frames[11][1][18] = 8'had;
frames[11][1][19] = 8'had;
frames[11][1][20] = 8'had;
frames[11][1][21] = 8'had;
frames[11][1][22] = 8'had;
frames[11][1][23] = 8'had;
frames[11][1][24] = 8'had;
frames[11][1][25] = 8'had;
frames[11][1][26] = 8'h89;
frames[11][1][27] = 8'h64;
frames[11][1][28] = 8'h40;
frames[11][1][29] = 8'h64;
frames[11][1][30] = 8'ha8;
frames[11][1][31] = 8'had;
frames[11][1][32] = 8'h8d;
frames[11][1][33] = 8'h44;
frames[11][1][34] = 8'h24;
frames[11][1][35] = 8'h24;
frames[11][1][36] = 8'h6d;
frames[11][1][37] = 8'hb6;
frames[11][1][38] = 8'hda;
frames[11][1][39] = 8'h6d;
frames[11][2][0] = 8'h00;
frames[11][2][1] = 8'h00;
frames[11][2][2] = 8'h00;
frames[11][2][3] = 8'h24;
frames[11][2][4] = 8'h49;
frames[11][2][5] = 8'h24;
frames[11][2][6] = 8'h20;
frames[11][2][7] = 8'h24;
frames[11][2][8] = 8'h44;
frames[11][2][9] = 8'h44;
frames[11][2][10] = 8'h64;
frames[11][2][11] = 8'h64;
frames[11][2][12] = 8'h89;
frames[11][2][13] = 8'had;
frames[11][2][14] = 8'had;
frames[11][2][15] = 8'had;
frames[11][2][16] = 8'had;
frames[11][2][17] = 8'had;
frames[11][2][18] = 8'had;
frames[11][2][19] = 8'had;
frames[11][2][20] = 8'had;
frames[11][2][21] = 8'had;
frames[11][2][22] = 8'had;
frames[11][2][23] = 8'had;
frames[11][2][24] = 8'had;
frames[11][2][25] = 8'had;
frames[11][2][26] = 8'had;
frames[11][2][27] = 8'h64;
frames[11][2][28] = 8'h40;
frames[11][2][29] = 8'h64;
frames[11][2][30] = 8'h64;
frames[11][2][31] = 8'h64;
frames[11][2][32] = 8'h24;
frames[11][2][33] = 8'h24;
frames[11][2][34] = 8'h24;
frames[11][2][35] = 8'h44;
frames[11][2][36] = 8'h92;
frames[11][2][37] = 8'h6d;
frames[11][2][38] = 8'h6d;
frames[11][2][39] = 8'h72;
frames[11][3][0] = 8'h00;
frames[11][3][1] = 8'h20;
frames[11][3][2] = 8'h44;
frames[11][3][3] = 8'h49;
frames[11][3][4] = 8'h49;
frames[11][3][5] = 8'h20;
frames[11][3][6] = 8'h20;
frames[11][3][7] = 8'h20;
frames[11][3][8] = 8'h24;
frames[11][3][9] = 8'h24;
frames[11][3][10] = 8'h24;
frames[11][3][11] = 8'h24;
frames[11][3][12] = 8'h24;
frames[11][3][13] = 8'h48;
frames[11][3][14] = 8'had;
frames[11][3][15] = 8'had;
frames[11][3][16] = 8'had;
frames[11][3][17] = 8'had;
frames[11][3][18] = 8'had;
frames[11][3][19] = 8'had;
frames[11][3][20] = 8'had;
frames[11][3][21] = 8'had;
frames[11][3][22] = 8'had;
frames[11][3][23] = 8'ha9;
frames[11][3][24] = 8'h89;
frames[11][3][25] = 8'h89;
frames[11][3][26] = 8'had;
frames[11][3][27] = 8'h89;
frames[11][3][28] = 8'h44;
frames[11][3][29] = 8'h40;
frames[11][3][30] = 8'h44;
frames[11][3][31] = 8'h44;
frames[11][3][32] = 8'h24;
frames[11][3][33] = 8'h24;
frames[11][3][34] = 8'h44;
frames[11][3][35] = 8'h68;
frames[11][3][36] = 8'h8d;
frames[11][3][37] = 8'h69;
frames[11][3][38] = 8'h48;
frames[11][3][39] = 8'h91;
frames[11][4][0] = 8'h24;
frames[11][4][1] = 8'h24;
frames[11][4][2] = 8'h44;
frames[11][4][3] = 8'h44;
frames[11][4][4] = 8'h24;
frames[11][4][5] = 8'h00;
frames[11][4][6] = 8'h00;
frames[11][4][7] = 8'h24;
frames[11][4][8] = 8'h24;
frames[11][4][9] = 8'h24;
frames[11][4][10] = 8'h20;
frames[11][4][11] = 8'h20;
frames[11][4][12] = 8'h20;
frames[11][4][13] = 8'h20;
frames[11][4][14] = 8'h68;
frames[11][4][15] = 8'had;
frames[11][4][16] = 8'had;
frames[11][4][17] = 8'had;
frames[11][4][18] = 8'had;
frames[11][4][19] = 8'had;
frames[11][4][20] = 8'had;
frames[11][4][21] = 8'had;
frames[11][4][22] = 8'h88;
frames[11][4][23] = 8'h88;
frames[11][4][24] = 8'h84;
frames[11][4][25] = 8'h88;
frames[11][4][26] = 8'h89;
frames[11][4][27] = 8'had;
frames[11][4][28] = 8'h89;
frames[11][4][29] = 8'h40;
frames[11][4][30] = 8'h44;
frames[11][4][31] = 8'h44;
frames[11][4][32] = 8'h44;
frames[11][4][33] = 8'h44;
frames[11][4][34] = 8'h44;
frames[11][4][35] = 8'h44;
frames[11][4][36] = 8'hb1;
frames[11][4][37] = 8'h8d;
frames[11][4][38] = 8'h8d;
frames[11][4][39] = 8'h8d;
frames[11][5][0] = 8'h24;
frames[11][5][1] = 8'h24;
frames[11][5][2] = 8'h44;
frames[11][5][3] = 8'h24;
frames[11][5][4] = 8'h00;
frames[11][5][5] = 8'h00;
frames[11][5][6] = 8'h00;
frames[11][5][7] = 8'h24;
frames[11][5][8] = 8'h24;
frames[11][5][9] = 8'h24;
frames[11][5][10] = 8'h20;
frames[11][5][11] = 8'h20;
frames[11][5][12] = 8'h20;
frames[11][5][13] = 8'h20;
frames[11][5][14] = 8'h44;
frames[11][5][15] = 8'had;
frames[11][5][16] = 8'had;
frames[11][5][17] = 8'had;
frames[11][5][18] = 8'had;
frames[11][5][19] = 8'had;
frames[11][5][20] = 8'had;
frames[11][5][21] = 8'h89;
frames[11][5][22] = 8'h89;
frames[11][5][23] = 8'h88;
frames[11][5][24] = 8'h64;
frames[11][5][25] = 8'h88;
frames[11][5][26] = 8'h88;
frames[11][5][27] = 8'ha9;
frames[11][5][28] = 8'had;
frames[11][5][29] = 8'h88;
frames[11][5][30] = 8'h64;
frames[11][5][31] = 8'h64;
frames[11][5][32] = 8'h64;
frames[11][5][33] = 8'h64;
frames[11][5][34] = 8'h64;
frames[11][5][35] = 8'h64;
frames[11][5][36] = 8'h68;
frames[11][5][37] = 8'hb1;
frames[11][5][38] = 8'hb1;
frames[11][5][39] = 8'h64;
frames[11][6][0] = 8'h24;
frames[11][6][1] = 8'h24;
frames[11][6][2] = 8'h44;
frames[11][6][3] = 8'h24;
frames[11][6][4] = 8'h24;
frames[11][6][5] = 8'h20;
frames[11][6][6] = 8'h44;
frames[11][6][7] = 8'h8d;
frames[11][6][8] = 8'h6d;
frames[11][6][9] = 8'h48;
frames[11][6][10] = 8'h24;
frames[11][6][11] = 8'h24;
frames[11][6][12] = 8'h24;
frames[11][6][13] = 8'h24;
frames[11][6][14] = 8'h20;
frames[11][6][15] = 8'h69;
frames[11][6][16] = 8'had;
frames[11][6][17] = 8'had;
frames[11][6][18] = 8'had;
frames[11][6][19] = 8'had;
frames[11][6][20] = 8'ha9;
frames[11][6][21] = 8'h88;
frames[11][6][22] = 8'h88;
frames[11][6][23] = 8'h89;
frames[11][6][24] = 8'h64;
frames[11][6][25] = 8'h64;
frames[11][6][26] = 8'h88;
frames[11][6][27] = 8'h89;
frames[11][6][28] = 8'had;
frames[11][6][29] = 8'had;
frames[11][6][30] = 8'h68;
frames[11][6][31] = 8'h64;
frames[11][6][32] = 8'h64;
frames[11][6][33] = 8'h64;
frames[11][6][34] = 8'h64;
frames[11][6][35] = 8'h64;
frames[11][6][36] = 8'h64;
frames[11][6][37] = 8'h64;
frames[11][6][38] = 8'h64;
frames[11][6][39] = 8'h68;
frames[11][7][0] = 8'h6d;
frames[11][7][1] = 8'h6d;
frames[11][7][2] = 8'h8d;
frames[11][7][3] = 8'h8d;
frames[11][7][4] = 8'h8d;
frames[11][7][5] = 8'h8d;
frames[11][7][6] = 8'h8d;
frames[11][7][7] = 8'h91;
frames[11][7][8] = 8'hb1;
frames[11][7][9] = 8'hb1;
frames[11][7][10] = 8'h8d;
frames[11][7][11] = 8'h68;
frames[11][7][12] = 8'h68;
frames[11][7][13] = 8'h68;
frames[11][7][14] = 8'h44;
frames[11][7][15] = 8'h48;
frames[11][7][16] = 8'had;
frames[11][7][17] = 8'had;
frames[11][7][18] = 8'had;
frames[11][7][19] = 8'had;
frames[11][7][20] = 8'h88;
frames[11][7][21] = 8'h84;
frames[11][7][22] = 8'h88;
frames[11][7][23] = 8'h89;
frames[11][7][24] = 8'had;
frames[11][7][25] = 8'h64;
frames[11][7][26] = 8'h64;
frames[11][7][27] = 8'h84;
frames[11][7][28] = 8'h89;
frames[11][7][29] = 8'had;
frames[11][7][30] = 8'h8d;
frames[11][7][31] = 8'h44;
frames[11][7][32] = 8'h44;
frames[11][7][33] = 8'h44;
frames[11][7][34] = 8'h64;
frames[11][7][35] = 8'h64;
frames[11][7][36] = 8'h64;
frames[11][7][37] = 8'h68;
frames[11][7][38] = 8'h68;
frames[11][7][39] = 8'h68;
frames[11][8][0] = 8'hb1;
frames[11][8][1] = 8'hb1;
frames[11][8][2] = 8'hb1;
frames[11][8][3] = 8'hb1;
frames[11][8][4] = 8'hb1;
frames[11][8][5] = 8'hb1;
frames[11][8][6] = 8'hb1;
frames[11][8][7] = 8'h91;
frames[11][8][8] = 8'hb1;
frames[11][8][9] = 8'hb1;
frames[11][8][10] = 8'h8d;
frames[11][8][11] = 8'h8d;
frames[11][8][12] = 8'h8d;
frames[11][8][13] = 8'h8d;
frames[11][8][14] = 8'h8d;
frames[11][8][15] = 8'h68;
frames[11][8][16] = 8'h89;
frames[11][8][17] = 8'had;
frames[11][8][18] = 8'had;
frames[11][8][19] = 8'h88;
frames[11][8][20] = 8'h64;
frames[11][8][21] = 8'h64;
frames[11][8][22] = 8'h84;
frames[11][8][23] = 8'h88;
frames[11][8][24] = 8'had;
frames[11][8][25] = 8'had;
frames[11][8][26] = 8'h44;
frames[11][8][27] = 8'h64;
frames[11][8][28] = 8'h84;
frames[11][8][29] = 8'ha9;
frames[11][8][30] = 8'had;
frames[11][8][31] = 8'h89;
frames[11][8][32] = 8'h44;
frames[11][8][33] = 8'h44;
frames[11][8][34] = 8'h44;
frames[11][8][35] = 8'h44;
frames[11][8][36] = 8'h44;
frames[11][8][37] = 8'h44;
frames[11][8][38] = 8'h44;
frames[11][8][39] = 8'h44;
frames[11][9][0] = 8'h8d;
frames[11][9][1] = 8'h8d;
frames[11][9][2] = 8'h88;
frames[11][9][3] = 8'h88;
frames[11][9][4] = 8'h8d;
frames[11][9][5] = 8'h8d;
frames[11][9][6] = 8'hb1;
frames[11][9][7] = 8'h88;
frames[11][9][8] = 8'h84;
frames[11][9][9] = 8'h64;
frames[11][9][10] = 8'h64;
frames[11][9][11] = 8'had;
frames[11][9][12] = 8'hb1;
frames[11][9][13] = 8'hb1;
frames[11][9][14] = 8'hb1;
frames[11][9][15] = 8'h91;
frames[11][9][16] = 8'h8d;
frames[11][9][17] = 8'h8d;
frames[11][9][18] = 8'had;
frames[11][9][19] = 8'h88;
frames[11][9][20] = 8'h64;
frames[11][9][21] = 8'h64;
frames[11][9][22] = 8'h64;
frames[11][9][23] = 8'h64;
frames[11][9][24] = 8'h89;
frames[11][9][25] = 8'had;
frames[11][9][26] = 8'h89;
frames[11][9][27] = 8'h44;
frames[11][9][28] = 8'h64;
frames[11][9][29] = 8'h88;
frames[11][9][30] = 8'had;
frames[11][9][31] = 8'hcd;
frames[11][9][32] = 8'h8d;
frames[11][9][33] = 8'h44;
frames[11][9][34] = 8'h24;
frames[11][9][35] = 8'h24;
frames[11][9][36] = 8'h24;
frames[11][9][37] = 8'h24;
frames[11][9][38] = 8'h24;
frames[11][9][39] = 8'h24;
frames[11][10][0] = 8'h8d;
frames[11][10][1] = 8'h88;
frames[11][10][2] = 8'h64;
frames[11][10][3] = 8'h88;
frames[11][10][4] = 8'hb1;
frames[11][10][5] = 8'hb1;
frames[11][10][6] = 8'ha8;
frames[11][10][7] = 8'h64;
frames[11][10][8] = 8'h84;
frames[11][10][9] = 8'h84;
frames[11][10][10] = 8'h64;
frames[11][10][11] = 8'hd1;
frames[11][10][12] = 8'hd6;
frames[11][10][13] = 8'hb5;
frames[11][10][14] = 8'hb1;
frames[11][10][15] = 8'hb2;
frames[11][10][16] = 8'hb1;
frames[11][10][17] = 8'h68;
frames[11][10][18] = 8'h88;
frames[11][10][19] = 8'h64;
frames[11][10][20] = 8'h64;
frames[11][10][21] = 8'h64;
frames[11][10][22] = 8'h64;
frames[11][10][23] = 8'h64;
frames[11][10][24] = 8'h88;
frames[11][10][25] = 8'h89;
frames[11][10][26] = 8'had;
frames[11][10][27] = 8'h88;
frames[11][10][28] = 8'h40;
frames[11][10][29] = 8'h64;
frames[11][10][30] = 8'ha9;
frames[11][10][31] = 8'hcd;
frames[11][10][32] = 8'had;
frames[11][10][33] = 8'h64;
frames[11][10][34] = 8'h24;
frames[11][10][35] = 8'h24;
frames[11][10][36] = 8'h24;
frames[11][10][37] = 8'h24;
frames[11][10][38] = 8'h24;
frames[11][10][39] = 8'h24;
frames[11][11][0] = 8'h88;
frames[11][11][1] = 8'h88;
frames[11][11][2] = 8'h84;
frames[11][11][3] = 8'h84;
frames[11][11][4] = 8'h88;
frames[11][11][5] = 8'hb1;
frames[11][11][6] = 8'had;
frames[11][11][7] = 8'h88;
frames[11][11][8] = 8'ha8;
frames[11][11][9] = 8'h84;
frames[11][11][10] = 8'h88;
frames[11][11][11] = 8'hd1;
frames[11][11][12] = 8'hd5;
frames[11][11][13] = 8'hd5;
frames[11][11][14] = 8'hd6;
frames[11][11][15] = 8'hd6;
frames[11][11][16] = 8'hb2;
frames[11][11][17] = 8'h44;
frames[11][11][18] = 8'h64;
frames[11][11][19] = 8'h44;
frames[11][11][20] = 8'h64;
frames[11][11][21] = 8'h64;
frames[11][11][22] = 8'h64;
frames[11][11][23] = 8'h64;
frames[11][11][24] = 8'h64;
frames[11][11][25] = 8'h88;
frames[11][11][26] = 8'h89;
frames[11][11][27] = 8'had;
frames[11][11][28] = 8'h89;
frames[11][11][29] = 8'h64;
frames[11][11][30] = 8'h84;
frames[11][11][31] = 8'ha9;
frames[11][11][32] = 8'had;
frames[11][11][33] = 8'h64;
frames[11][11][34] = 8'h24;
frames[11][11][35] = 8'h24;
frames[11][11][36] = 8'h24;
frames[11][11][37] = 8'h24;
frames[11][11][38] = 8'h24;
frames[11][11][39] = 8'h24;
frames[11][12][0] = 8'hcd;
frames[11][12][1] = 8'h84;
frames[11][12][2] = 8'h84;
frames[11][12][3] = 8'h80;
frames[11][12][4] = 8'h88;
frames[11][12][5] = 8'hcd;
frames[11][12][6] = 8'hb1;
frames[11][12][7] = 8'hb1;
frames[11][12][8] = 8'had;
frames[11][12][9] = 8'h88;
frames[11][12][10] = 8'h84;
frames[11][12][11] = 8'ha8;
frames[11][12][12] = 8'h8d;
frames[11][12][13] = 8'hd1;
frames[11][12][14] = 8'hd6;
frames[11][12][15] = 8'hd6;
frames[11][12][16] = 8'h91;
frames[11][12][17] = 8'h44;
frames[11][12][18] = 8'h44;
frames[11][12][19] = 8'h44;
frames[11][12][20] = 8'h44;
frames[11][12][21] = 8'h44;
frames[11][12][22] = 8'h64;
frames[11][12][23] = 8'h64;
frames[11][12][24] = 8'h64;
frames[11][12][25] = 8'h64;
frames[11][12][26] = 8'h88;
frames[11][12][27] = 8'h89;
frames[11][12][28] = 8'had;
frames[11][12][29] = 8'had;
frames[11][12][30] = 8'h84;
frames[11][12][31] = 8'h88;
frames[11][12][32] = 8'ha8;
frames[11][12][33] = 8'h84;
frames[11][12][34] = 8'h44;
frames[11][12][35] = 8'h40;
frames[11][12][36] = 8'h24;
frames[11][12][37] = 8'h24;
frames[11][12][38] = 8'h24;
frames[11][12][39] = 8'h24;
frames[11][13][0] = 8'hf6;
frames[11][13][1] = 8'had;
frames[11][13][2] = 8'ha4;
frames[11][13][3] = 8'h84;
frames[11][13][4] = 8'h84;
frames[11][13][5] = 8'ha8;
frames[11][13][6] = 8'h88;
frames[11][13][7] = 8'had;
frames[11][13][8] = 8'hd5;
frames[11][13][9] = 8'hb1;
frames[11][13][10] = 8'hd1;
frames[11][13][11] = 8'had;
frames[11][13][12] = 8'h88;
frames[11][13][13] = 8'hd1;
frames[11][13][14] = 8'hb1;
frames[11][13][15] = 8'hb5;
frames[11][13][16] = 8'h69;
frames[11][13][17] = 8'h44;
frames[11][13][18] = 8'h44;
frames[11][13][19] = 8'h44;
frames[11][13][20] = 8'h44;
frames[11][13][21] = 8'h48;
frames[11][13][22] = 8'h44;
frames[11][13][23] = 8'h44;
frames[11][13][24] = 8'h64;
frames[11][13][25] = 8'h64;
frames[11][13][26] = 8'h64;
frames[11][13][27] = 8'h68;
frames[11][13][28] = 8'had;
frames[11][13][29] = 8'had;
frames[11][13][30] = 8'h88;
frames[11][13][31] = 8'h64;
frames[11][13][32] = 8'h84;
frames[11][13][33] = 8'h80;
frames[11][13][34] = 8'h44;
frames[11][13][35] = 8'h40;
frames[11][13][36] = 8'h24;
frames[11][13][37] = 8'h24;
frames[11][13][38] = 8'h24;
frames[11][13][39] = 8'h24;
frames[11][14][0] = 8'hd1;
frames[11][14][1] = 8'hd5;
frames[11][14][2] = 8'hac;
frames[11][14][3] = 8'h64;
frames[11][14][4] = 8'h84;
frames[11][14][5] = 8'h84;
frames[11][14][6] = 8'h88;
frames[11][14][7] = 8'hcd;
frames[11][14][8] = 8'hb1;
frames[11][14][9] = 8'hb1;
frames[11][14][10] = 8'hd6;
frames[11][14][11] = 8'hda;
frames[11][14][12] = 8'hb5;
frames[11][14][13] = 8'hb1;
frames[11][14][14] = 8'hb6;
frames[11][14][15] = 8'h6d;
frames[11][14][16] = 8'h44;
frames[11][14][17] = 8'h44;
frames[11][14][18] = 8'h44;
frames[11][14][19] = 8'h44;
frames[11][14][20] = 8'h48;
frames[11][14][21] = 8'h44;
frames[11][14][22] = 8'h48;
frames[11][14][23] = 8'h69;
frames[11][14][24] = 8'h68;
frames[11][14][25] = 8'h64;
frames[11][14][26] = 8'h64;
frames[11][14][27] = 8'h89;
frames[11][14][28] = 8'h88;
frames[11][14][29] = 8'h8d;
frames[11][14][30] = 8'h88;
frames[11][14][31] = 8'h64;
frames[11][14][32] = 8'h60;
frames[11][14][33] = 8'h60;
frames[11][14][34] = 8'h64;
frames[11][14][35] = 8'h44;
frames[11][14][36] = 8'h24;
frames[11][14][37] = 8'h24;
frames[11][14][38] = 8'h24;
frames[11][14][39] = 8'h24;
frames[11][15][0] = 8'h88;
frames[11][15][1] = 8'hb1;
frames[11][15][2] = 8'hd1;
frames[11][15][3] = 8'hac;
frames[11][15][4] = 8'h88;
frames[11][15][5] = 8'ha8;
frames[11][15][6] = 8'h8c;
frames[11][15][7] = 8'hb1;
frames[11][15][8] = 8'hd5;
frames[11][15][9] = 8'hd5;
frames[11][15][10] = 8'hd5;
frames[11][15][11] = 8'hd5;
frames[11][15][12] = 8'hb1;
frames[11][15][13] = 8'h91;
frames[11][15][14] = 8'h69;
frames[11][15][15] = 8'h24;
frames[11][15][16] = 8'h24;
frames[11][15][17] = 8'h44;
frames[11][15][18] = 8'h44;
frames[11][15][19] = 8'h6d;
frames[11][15][20] = 8'hb1;
frames[11][15][21] = 8'h88;
frames[11][15][22] = 8'h88;
frames[11][15][23] = 8'h8c;
frames[11][15][24] = 8'h8d;
frames[11][15][25] = 8'had;
frames[11][15][26] = 8'h8d;
frames[11][15][27] = 8'h8d;
frames[11][15][28] = 8'had;
frames[11][15][29] = 8'hb1;
frames[11][15][30] = 8'h8c;
frames[11][15][31] = 8'h88;
frames[11][15][32] = 8'h64;
frames[11][15][33] = 8'h64;
frames[11][15][34] = 8'h64;
frames[11][15][35] = 8'h64;
frames[11][15][36] = 8'h48;
frames[11][15][37] = 8'h6d;
frames[11][15][38] = 8'h24;
frames[11][15][39] = 8'h24;
frames[11][16][0] = 8'h8d;
frames[11][16][1] = 8'hd6;
frames[11][16][2] = 8'hd6;
frames[11][16][3] = 8'hd6;
frames[11][16][4] = 8'hb1;
frames[11][16][5] = 8'h8d;
frames[11][16][6] = 8'had;
frames[11][16][7] = 8'hd5;
frames[11][16][8] = 8'hb5;
frames[11][16][9] = 8'hd5;
frames[11][16][10] = 8'hb5;
frames[11][16][11] = 8'hb1;
frames[11][16][12] = 8'h68;
frames[11][16][13] = 8'h44;
frames[11][16][14] = 8'h24;
frames[11][16][15] = 8'h44;
frames[11][16][16] = 8'h48;
frames[11][16][17] = 8'h69;
frames[11][16][18] = 8'h8d;
frames[11][16][19] = 8'had;
frames[11][16][20] = 8'hb1;
frames[11][16][21] = 8'hd1;
frames[11][16][22] = 8'had;
frames[11][16][23] = 8'hac;
frames[11][16][24] = 8'h8c;
frames[11][16][25] = 8'hd1;
frames[11][16][26] = 8'hd5;
frames[11][16][27] = 8'hb1;
frames[11][16][28] = 8'hb1;
frames[11][16][29] = 8'hb1;
frames[11][16][30] = 8'hb1;
frames[11][16][31] = 8'hb1;
frames[11][16][32] = 8'hb1;
frames[11][16][33] = 8'h8c;
frames[11][16][34] = 8'had;
frames[11][16][35] = 8'hd1;
frames[11][16][36] = 8'hb1;
frames[11][16][37] = 8'hb1;
frames[11][16][38] = 8'h48;
frames[11][16][39] = 8'h44;
frames[11][17][0] = 8'hd6;
frames[11][17][1] = 8'hd6;
frames[11][17][2] = 8'hd5;
frames[11][17][3] = 8'hb5;
frames[11][17][4] = 8'hd6;
frames[11][17][5] = 8'hb1;
frames[11][17][6] = 8'hb5;
frames[11][17][7] = 8'hd5;
frames[11][17][8] = 8'hd6;
frames[11][17][9] = 8'h91;
frames[11][17][10] = 8'h48;
frames[11][17][11] = 8'h20;
frames[11][17][12] = 8'h20;
frames[11][17][13] = 8'h20;
frames[11][17][14] = 8'h48;
frames[11][17][15] = 8'h8d;
frames[11][17][16] = 8'h88;
frames[11][17][17] = 8'h88;
frames[11][17][18] = 8'h88;
frames[11][17][19] = 8'ha8;
frames[11][17][20] = 8'hb1;
frames[11][17][21] = 8'hd1;
frames[11][17][22] = 8'had;
frames[11][17][23] = 8'hb1;
frames[11][17][24] = 8'hd5;
frames[11][17][25] = 8'hd6;
frames[11][17][26] = 8'hd6;
frames[11][17][27] = 8'hb1;
frames[11][17][28] = 8'hb1;
frames[11][17][29] = 8'hb1;
frames[11][17][30] = 8'hb1;
frames[11][17][31] = 8'hd6;
frames[11][17][32] = 8'hd5;
frames[11][17][33] = 8'hb1;
frames[11][17][34] = 8'hd6;
frames[11][17][35] = 8'hd6;
frames[11][17][36] = 8'hb5;
frames[11][17][37] = 8'hb5;
frames[11][17][38] = 8'h91;
frames[11][17][39] = 8'h6d;
frames[11][18][0] = 8'hda;
frames[11][18][1] = 8'hd6;
frames[11][18][2] = 8'hd6;
frames[11][18][3] = 8'hd6;
frames[11][18][4] = 8'hd6;
frames[11][18][5] = 8'hb1;
frames[11][18][6] = 8'h91;
frames[11][18][7] = 8'h6c;
frames[11][18][8] = 8'h44;
frames[11][18][9] = 8'h20;
frames[11][18][10] = 8'h20;
frames[11][18][11] = 8'h20;
frames[11][18][12] = 8'h20;
frames[11][18][13] = 8'h48;
frames[11][18][14] = 8'hb1;
frames[11][18][15] = 8'hb1;
frames[11][18][16] = 8'hcd;
frames[11][18][17] = 8'ha8;
frames[11][18][18] = 8'ha4;
frames[11][18][19] = 8'ha4;
frames[11][18][20] = 8'hd1;
frames[11][18][21] = 8'hd1;
frames[11][18][22] = 8'hb1;
frames[11][18][23] = 8'hb1;
frames[11][18][24] = 8'hd5;
frames[11][18][25] = 8'hd6;
frames[11][18][26] = 8'hd6;
frames[11][18][27] = 8'hd5;
frames[11][18][28] = 8'hda;
frames[11][18][29] = 8'hd5;
frames[11][18][30] = 8'hb1;
frames[11][18][31] = 8'hd5;
frames[11][18][32] = 8'hd5;
frames[11][18][33] = 8'hd1;
frames[11][18][34] = 8'hd6;
frames[11][18][35] = 8'hd6;
frames[11][18][36] = 8'hd6;
frames[11][18][37] = 8'hb1;
frames[11][18][38] = 8'hb1;
frames[11][18][39] = 8'h91;
frames[11][19][0] = 8'h6d;
frames[11][19][1] = 8'h8d;
frames[11][19][2] = 8'h8d;
frames[11][19][3] = 8'h6d;
frames[11][19][4] = 8'h48;
frames[11][19][5] = 8'h44;
frames[11][19][6] = 8'h24;
frames[11][19][7] = 8'h24;
frames[11][19][8] = 8'h24;
frames[11][19][9] = 8'h24;
frames[11][19][10] = 8'h24;
frames[11][19][11] = 8'h24;
frames[11][19][12] = 8'h69;
frames[11][19][13] = 8'hb1;
frames[11][19][14] = 8'hd6;
frames[11][19][15] = 8'hda;
frames[11][19][16] = 8'hd1;
frames[11][19][17] = 8'h88;
frames[11][19][18] = 8'h84;
frames[11][19][19] = 8'h84;
frames[11][19][20] = 8'had;
frames[11][19][21] = 8'hd1;
frames[11][19][22] = 8'had;
frames[11][19][23] = 8'had;
frames[11][19][24] = 8'hd5;
frames[11][19][25] = 8'hd6;
frames[11][19][26] = 8'hd6;
frames[11][19][27] = 8'hb1;
frames[11][19][28] = 8'hd6;
frames[11][19][29] = 8'hd5;
frames[11][19][30] = 8'ha8;
frames[11][19][31] = 8'h88;
frames[11][19][32] = 8'h84;
frames[11][19][33] = 8'ha4;
frames[11][19][34] = 8'had;
frames[11][19][35] = 8'hd6;
frames[11][19][36] = 8'hd6;
frames[11][19][37] = 8'hb1;
frames[11][19][38] = 8'hb1;
frames[11][19][39] = 8'h91;
frames[11][20][0] = 8'h24;
frames[11][20][1] = 8'h24;
frames[11][20][2] = 8'h24;
frames[11][20][3] = 8'h24;
frames[11][20][4] = 8'h24;
frames[11][20][5] = 8'h24;
frames[11][20][6] = 8'h24;
frames[11][20][7] = 8'h24;
frames[11][20][8] = 8'h24;
frames[11][20][9] = 8'h24;
frames[11][20][10] = 8'h24;
frames[11][20][11] = 8'h44;
frames[11][20][12] = 8'h91;
frames[11][20][13] = 8'hb1;
frames[11][20][14] = 8'hd6;
frames[11][20][15] = 8'hd1;
frames[11][20][16] = 8'ha4;
frames[11][20][17] = 8'ha4;
frames[11][20][18] = 8'ha4;
frames[11][20][19] = 8'ha4;
frames[11][20][20] = 8'had;
frames[11][20][21] = 8'hb1;
frames[11][20][22] = 8'hcd;
frames[11][20][23] = 8'ha8;
frames[11][20][24] = 8'ha8;
frames[11][20][25] = 8'hcd;
frames[11][20][26] = 8'hd1;
frames[11][20][27] = 8'hb1;
frames[11][20][28] = 8'hd5;
frames[11][20][29] = 8'hb1;
frames[11][20][30] = 8'h84;
frames[11][20][31] = 8'ha4;
frames[11][20][32] = 8'h84;
frames[11][20][33] = 8'ha4;
frames[11][20][34] = 8'h88;
frames[11][20][35] = 8'hd1;
frames[11][20][36] = 8'hd6;
frames[11][20][37] = 8'hd6;
frames[11][20][38] = 8'hb1;
frames[11][20][39] = 8'hb1;
frames[11][21][0] = 8'h48;
frames[11][21][1] = 8'h44;
frames[11][21][2] = 8'h24;
frames[11][21][3] = 8'h24;
frames[11][21][4] = 8'h24;
frames[11][21][5] = 8'h24;
frames[11][21][6] = 8'h24;
frames[11][21][7] = 8'h24;
frames[11][21][8] = 8'h24;
frames[11][21][9] = 8'h24;
frames[11][21][10] = 8'h24;
frames[11][21][11] = 8'h24;
frames[11][21][12] = 8'h91;
frames[11][21][13] = 8'h91;
frames[11][21][14] = 8'hd1;
frames[11][21][15] = 8'hb1;
frames[11][21][16] = 8'ha8;
frames[11][21][17] = 8'ha8;
frames[11][21][18] = 8'hcd;
frames[11][21][19] = 8'hd1;
frames[11][21][20] = 8'hb1;
frames[11][21][21] = 8'h8d;
frames[11][21][22] = 8'hd1;
frames[11][21][23] = 8'hd1;
frames[11][21][24] = 8'hc8;
frames[11][21][25] = 8'ha8;
frames[11][21][26] = 8'ha8;
frames[11][21][27] = 8'ha8;
frames[11][21][28] = 8'hb1;
frames[11][21][29] = 8'hb1;
frames[11][21][30] = 8'ha4;
frames[11][21][31] = 8'h84;
frames[11][21][32] = 8'h84;
frames[11][21][33] = 8'ha4;
frames[11][21][34] = 8'had;
frames[11][21][35] = 8'hd1;
frames[11][21][36] = 8'hb1;
frames[11][21][37] = 8'hb1;
frames[11][21][38] = 8'h91;
frames[11][21][39] = 8'h68;
frames[11][22][0] = 8'h49;
frames[11][22][1] = 8'h48;
frames[11][22][2] = 8'h48;
frames[11][22][3] = 8'h44;
frames[11][22][4] = 8'h24;
frames[11][22][5] = 8'h24;
frames[11][22][6] = 8'h24;
frames[11][22][7] = 8'h24;
frames[11][22][8] = 8'h24;
frames[11][22][9] = 8'h24;
frames[11][22][10] = 8'h24;
frames[11][22][11] = 8'h24;
frames[11][22][12] = 8'h69;
frames[11][22][13] = 8'hb1;
frames[11][22][14] = 8'hb1;
frames[11][22][15] = 8'hb1;
frames[11][22][16] = 8'hd5;
frames[11][22][17] = 8'hd1;
frames[11][22][18] = 8'had;
frames[11][22][19] = 8'hd5;
frames[11][22][20] = 8'hb5;
frames[11][22][21] = 8'hb1;
frames[11][22][22] = 8'hd5;
frames[11][22][23] = 8'hb1;
frames[11][22][24] = 8'hd1;
frames[11][22][25] = 8'hac;
frames[11][22][26] = 8'ha8;
frames[11][22][27] = 8'hac;
frames[11][22][28] = 8'hb1;
frames[11][22][29] = 8'hb1;
frames[11][22][30] = 8'had;
frames[11][22][31] = 8'hac;
frames[11][22][32] = 8'hac;
frames[11][22][33] = 8'hd1;
frames[11][22][34] = 8'hd6;
frames[11][22][35] = 8'hb1;
frames[11][22][36] = 8'hb6;
frames[11][22][37] = 8'h8d;
frames[11][22][38] = 8'h24;
frames[11][22][39] = 8'h24;
frames[11][23][0] = 8'h44;
frames[11][23][1] = 8'h48;
frames[11][23][2] = 8'h48;
frames[11][23][3] = 8'h69;
frames[11][23][4] = 8'h49;
frames[11][23][5] = 8'h48;
frames[11][23][6] = 8'h44;
frames[11][23][7] = 8'h24;
frames[11][23][8] = 8'h24;
frames[11][23][9] = 8'h24;
frames[11][23][10] = 8'h24;
frames[11][23][11] = 8'h24;
frames[11][23][12] = 8'h24;
frames[11][23][13] = 8'h6d;
frames[11][23][14] = 8'hb1;
frames[11][23][15] = 8'hb2;
frames[11][23][16] = 8'hd6;
frames[11][23][17] = 8'hd6;
frames[11][23][18] = 8'hd6;
frames[11][23][19] = 8'hd6;
frames[11][23][20] = 8'hd5;
frames[11][23][21] = 8'hd5;
frames[11][23][22] = 8'hd6;
frames[11][23][23] = 8'hd5;
frames[11][23][24] = 8'hd6;
frames[11][23][25] = 8'hd6;
frames[11][23][26] = 8'hd6;
frames[11][23][27] = 8'hd6;
frames[11][23][28] = 8'hd5;
frames[11][23][29] = 8'hd5;
frames[11][23][30] = 8'hfa;
frames[11][23][31] = 8'hd6;
frames[11][23][32] = 8'hd5;
frames[11][23][33] = 8'hb1;
frames[11][23][34] = 8'hb1;
frames[11][23][35] = 8'h6d;
frames[11][23][36] = 8'h44;
frames[11][23][37] = 8'h24;
frames[11][23][38] = 8'h44;
frames[11][23][39] = 8'h48;
frames[11][24][0] = 8'h68;
frames[11][24][1] = 8'h48;
frames[11][24][2] = 8'h44;
frames[11][24][3] = 8'h44;
frames[11][24][4] = 8'h44;
frames[11][24][5] = 8'h44;
frames[11][24][6] = 8'h49;
frames[11][24][7] = 8'h49;
frames[11][24][8] = 8'h48;
frames[11][24][9] = 8'h44;
frames[11][24][10] = 8'h24;
frames[11][24][11] = 8'h24;
frames[11][24][12] = 8'h24;
frames[11][24][13] = 8'h24;
frames[11][24][14] = 8'h44;
frames[11][24][15] = 8'h6d;
frames[11][24][16] = 8'hb1;
frames[11][24][17] = 8'hd6;
frames[11][24][18] = 8'hd6;
frames[11][24][19] = 8'hd6;
frames[11][24][20] = 8'hd6;
frames[11][24][21] = 8'hd5;
frames[11][24][22] = 8'hb5;
frames[11][24][23] = 8'hd6;
frames[11][24][24] = 8'hd6;
frames[11][24][25] = 8'hd6;
frames[11][24][26] = 8'hd6;
frames[11][24][27] = 8'hd6;
frames[11][24][28] = 8'hd6;
frames[11][24][29] = 8'hb6;
frames[11][24][30] = 8'hb1;
frames[11][24][31] = 8'h8d;
frames[11][24][32] = 8'h6d;
frames[11][24][33] = 8'h44;
frames[11][24][34] = 8'h20;
frames[11][24][35] = 8'h20;
frames[11][24][36] = 8'h24;
frames[11][24][37] = 8'h44;
frames[11][24][38] = 8'h48;
frames[11][24][39] = 8'h49;
frames[11][25][0] = 8'h8d;
frames[11][25][1] = 8'h8d;
frames[11][25][2] = 8'h8d;
frames[11][25][3] = 8'h68;
frames[11][25][4] = 8'h68;
frames[11][25][5] = 8'h44;
frames[11][25][6] = 8'h44;
frames[11][25][7] = 8'h44;
frames[11][25][8] = 8'h44;
frames[11][25][9] = 8'h44;
frames[11][25][10] = 8'h48;
frames[11][25][11] = 8'h48;
frames[11][25][12] = 8'h48;
frames[11][25][13] = 8'h44;
frames[11][25][14] = 8'h24;
frames[11][25][15] = 8'h24;
frames[11][25][16] = 8'h24;
frames[11][25][17] = 8'h24;
frames[11][25][18] = 8'h44;
frames[11][25][19] = 8'h48;
frames[11][25][20] = 8'h68;
frames[11][25][21] = 8'h68;
frames[11][25][22] = 8'h68;
frames[11][25][23] = 8'h48;
frames[11][25][24] = 8'h68;
frames[11][25][25] = 8'h68;
frames[11][25][26] = 8'h48;
frames[11][25][27] = 8'h44;
frames[11][25][28] = 8'h44;
frames[11][25][29] = 8'h44;
frames[11][25][30] = 8'h24;
frames[11][25][31] = 8'h20;
frames[11][25][32] = 8'h00;
frames[11][25][33] = 8'h00;
frames[11][25][34] = 8'h24;
frames[11][25][35] = 8'h44;
frames[11][25][36] = 8'h49;
frames[11][25][37] = 8'h49;
frames[11][25][38] = 8'h48;
frames[11][25][39] = 8'h48;
frames[11][26][0] = 8'hb1;
frames[11][26][1] = 8'hb1;
frames[11][26][2] = 8'hb1;
frames[11][26][3] = 8'had;
frames[11][26][4] = 8'h8c;
frames[11][26][5] = 8'h8c;
frames[11][26][6] = 8'h68;
frames[11][26][7] = 8'h64;
frames[11][26][8] = 8'h44;
frames[11][26][9] = 8'h44;
frames[11][26][10] = 8'h44;
frames[11][26][11] = 8'h44;
frames[11][26][12] = 8'h44;
frames[11][26][13] = 8'h48;
frames[11][26][14] = 8'h48;
frames[11][26][15] = 8'h48;
frames[11][26][16] = 8'h44;
frames[11][26][17] = 8'h24;
frames[11][26][18] = 8'h20;
frames[11][26][19] = 8'h00;
frames[11][26][20] = 8'h00;
frames[11][26][21] = 8'h00;
frames[11][26][22] = 8'h00;
frames[11][26][23] = 8'h00;
frames[11][26][24] = 8'h00;
frames[11][26][25] = 8'h00;
frames[11][26][26] = 8'h00;
frames[11][26][27] = 8'h00;
frames[11][26][28] = 8'h00;
frames[11][26][29] = 8'h00;
frames[11][26][30] = 8'h00;
frames[11][26][31] = 8'h00;
frames[11][26][32] = 8'h20;
frames[11][26][33] = 8'h24;
frames[11][26][34] = 8'h44;
frames[11][26][35] = 8'h49;
frames[11][26][36] = 8'h68;
frames[11][26][37] = 8'h48;
frames[11][26][38] = 8'h44;
frames[11][26][39] = 8'h44;
frames[11][27][0] = 8'hb1;
frames[11][27][1] = 8'hb1;
frames[11][27][2] = 8'hb1;
frames[11][27][3] = 8'hb1;
frames[11][27][4] = 8'hb1;
frames[11][27][5] = 8'had;
frames[11][27][6] = 8'had;
frames[11][27][7] = 8'h8c;
frames[11][27][8] = 8'h88;
frames[11][27][9] = 8'h68;
frames[11][27][10] = 8'h44;
frames[11][27][11] = 8'h44;
frames[11][27][12] = 8'h44;
frames[11][27][13] = 8'h44;
frames[11][27][14] = 8'h44;
frames[11][27][15] = 8'h44;
frames[11][27][16] = 8'h48;
frames[11][27][17] = 8'h48;
frames[11][27][18] = 8'h48;
frames[11][27][19] = 8'h44;
frames[11][27][20] = 8'h44;
frames[11][27][21] = 8'h24;
frames[11][27][22] = 8'h24;
frames[11][27][23] = 8'h24;
frames[11][27][24] = 8'h24;
frames[11][27][25] = 8'h24;
frames[11][27][26] = 8'h24;
frames[11][27][27] = 8'h24;
frames[11][27][28] = 8'h24;
frames[11][27][29] = 8'h24;
frames[11][27][30] = 8'h24;
frames[11][27][31] = 8'h24;
frames[11][27][32] = 8'h44;
frames[11][27][33] = 8'h49;
frames[11][27][34] = 8'h69;
frames[11][27][35] = 8'h69;
frames[11][27][36] = 8'h44;
frames[11][27][37] = 8'h44;
frames[11][27][38] = 8'h44;
frames[11][27][39] = 8'h44;
frames[11][28][0] = 8'hb1;
frames[11][28][1] = 8'hb1;
frames[11][28][2] = 8'hb1;
frames[11][28][3] = 8'hb1;
frames[11][28][4] = 8'hb1;
frames[11][28][5] = 8'hb1;
frames[11][28][6] = 8'hb1;
frames[11][28][7] = 8'had;
frames[11][28][8] = 8'had;
frames[11][28][9] = 8'hac;
frames[11][28][10] = 8'h8c;
frames[11][28][11] = 8'h8c;
frames[11][28][12] = 8'h68;
frames[11][28][13] = 8'h68;
frames[11][28][14] = 8'h44;
frames[11][28][15] = 8'h44;
frames[11][28][16] = 8'h44;
frames[11][28][17] = 8'h44;
frames[11][28][18] = 8'h44;
frames[11][28][19] = 8'h44;
frames[11][28][20] = 8'h48;
frames[11][28][21] = 8'h48;
frames[11][28][22] = 8'h44;
frames[11][28][23] = 8'h44;
frames[11][28][24] = 8'h44;
frames[11][28][25] = 8'h44;
frames[11][28][26] = 8'h24;
frames[11][28][27] = 8'h24;
frames[11][28][28] = 8'h24;
frames[11][28][29] = 8'h24;
frames[11][28][30] = 8'h44;
frames[11][28][31] = 8'h48;
frames[11][28][32] = 8'h69;
frames[11][28][33] = 8'h69;
frames[11][28][34] = 8'h44;
frames[11][28][35] = 8'h44;
frames[11][28][36] = 8'h44;
frames[11][28][37] = 8'h44;
frames[11][28][38] = 8'h44;
frames[11][28][39] = 8'h44;
frames[11][29][0] = 8'hb1;
frames[11][29][1] = 8'hb1;
frames[11][29][2] = 8'hb1;
frames[11][29][3] = 8'hb1;
frames[11][29][4] = 8'hb1;
frames[11][29][5] = 8'hb1;
frames[11][29][6] = 8'hb1;
frames[11][29][7] = 8'had;
frames[11][29][8] = 8'had;
frames[11][29][9] = 8'had;
frames[11][29][10] = 8'had;
frames[11][29][11] = 8'had;
frames[11][29][12] = 8'h8d;
frames[11][29][13] = 8'h8c;
frames[11][29][14] = 8'h88;
frames[11][29][15] = 8'h68;
frames[11][29][16] = 8'h48;
frames[11][29][17] = 8'h44;
frames[11][29][18] = 8'h44;
frames[11][29][19] = 8'h44;
frames[11][29][20] = 8'h44;
frames[11][29][21] = 8'h44;
frames[11][29][22] = 8'h44;
frames[11][29][23] = 8'h48;
frames[11][29][24] = 8'h68;
frames[11][29][25] = 8'h48;
frames[11][29][26] = 8'h44;
frames[11][29][27] = 8'h44;
frames[11][29][28] = 8'h44;
frames[11][29][29] = 8'h48;
frames[11][29][30] = 8'h69;
frames[11][29][31] = 8'h48;
frames[11][29][32] = 8'h44;
frames[11][29][33] = 8'h44;
frames[11][29][34] = 8'h44;
frames[11][29][35] = 8'h44;
frames[11][29][36] = 8'h44;
frames[11][29][37] = 8'h44;
frames[11][29][38] = 8'h44;
frames[11][29][39] = 8'h44;
frames[12][0][0] = 8'h68;
frames[12][0][1] = 8'h68;
frames[12][0][2] = 8'h88;
frames[12][0][3] = 8'h88;
frames[12][0][4] = 8'h88;
frames[12][0][5] = 8'h88;
frames[12][0][6] = 8'h89;
frames[12][0][7] = 8'h89;
frames[12][0][8] = 8'ha9;
frames[12][0][9] = 8'ha9;
frames[12][0][10] = 8'ha9;
frames[12][0][11] = 8'had;
frames[12][0][12] = 8'had;
frames[12][0][13] = 8'had;
frames[12][0][14] = 8'had;
frames[12][0][15] = 8'had;
frames[12][0][16] = 8'had;
frames[12][0][17] = 8'had;
frames[12][0][18] = 8'h88;
frames[12][0][19] = 8'h88;
frames[12][0][20] = 8'h88;
frames[12][0][21] = 8'had;
frames[12][0][22] = 8'had;
frames[12][0][23] = 8'h64;
frames[12][0][24] = 8'h89;
frames[12][0][25] = 8'ha9;
frames[12][0][26] = 8'h89;
frames[12][0][27] = 8'h40;
frames[12][0][28] = 8'h60;
frames[12][0][29] = 8'h40;
frames[12][0][30] = 8'h84;
frames[12][0][31] = 8'h88;
frames[12][0][32] = 8'h8d;
frames[12][0][33] = 8'had;
frames[12][0][34] = 8'h24;
frames[12][0][35] = 8'h24;
frames[12][0][36] = 8'h24;
frames[12][0][37] = 8'h6d;
frames[12][0][38] = 8'h6d;
frames[12][0][39] = 8'h69;
frames[12][1][0] = 8'h68;
frames[12][1][1] = 8'h68;
frames[12][1][2] = 8'h68;
frames[12][1][3] = 8'h88;
frames[12][1][4] = 8'h88;
frames[12][1][5] = 8'h88;
frames[12][1][6] = 8'h89;
frames[12][1][7] = 8'h89;
frames[12][1][8] = 8'h89;
frames[12][1][9] = 8'h89;
frames[12][1][10] = 8'had;
frames[12][1][11] = 8'had;
frames[12][1][12] = 8'had;
frames[12][1][13] = 8'had;
frames[12][1][14] = 8'had;
frames[12][1][15] = 8'had;
frames[12][1][16] = 8'had;
frames[12][1][17] = 8'had;
frames[12][1][18] = 8'h88;
frames[12][1][19] = 8'h64;
frames[12][1][20] = 8'h88;
frames[12][1][21] = 8'h89;
frames[12][1][22] = 8'had;
frames[12][1][23] = 8'h88;
frames[12][1][24] = 8'h84;
frames[12][1][25] = 8'ha9;
frames[12][1][26] = 8'had;
frames[12][1][27] = 8'h64;
frames[12][1][28] = 8'h60;
frames[12][1][29] = 8'h60;
frames[12][1][30] = 8'h60;
frames[12][1][31] = 8'h84;
frames[12][1][32] = 8'hb1;
frames[12][1][33] = 8'h8d;
frames[12][1][34] = 8'h24;
frames[12][1][35] = 8'h24;
frames[12][1][36] = 8'h6d;
frames[12][1][37] = 8'hb6;
frames[12][1][38] = 8'hda;
frames[12][1][39] = 8'h6d;
frames[12][2][0] = 8'h44;
frames[12][2][1] = 8'h44;
frames[12][2][2] = 8'h68;
frames[12][2][3] = 8'h88;
frames[12][2][4] = 8'h88;
frames[12][2][5] = 8'h89;
frames[12][2][6] = 8'h89;
frames[12][2][7] = 8'h89;
frames[12][2][8] = 8'h88;
frames[12][2][9] = 8'h89;
frames[12][2][10] = 8'had;
frames[12][2][11] = 8'had;
frames[12][2][12] = 8'had;
frames[12][2][13] = 8'had;
frames[12][2][14] = 8'had;
frames[12][2][15] = 8'had;
frames[12][2][16] = 8'had;
frames[12][2][17] = 8'had;
frames[12][2][18] = 8'ha9;
frames[12][2][19] = 8'h64;
frames[12][2][20] = 8'h64;
frames[12][2][21] = 8'h88;
frames[12][2][22] = 8'had;
frames[12][2][23] = 8'had;
frames[12][2][24] = 8'h84;
frames[12][2][25] = 8'h89;
frames[12][2][26] = 8'had;
frames[12][2][27] = 8'ha9;
frames[12][2][28] = 8'h60;
frames[12][2][29] = 8'h60;
frames[12][2][30] = 8'h84;
frames[12][2][31] = 8'ha9;
frames[12][2][32] = 8'h8d;
frames[12][2][33] = 8'h44;
frames[12][2][34] = 8'h24;
frames[12][2][35] = 8'h44;
frames[12][2][36] = 8'h92;
frames[12][2][37] = 8'h69;
frames[12][2][38] = 8'h6d;
frames[12][2][39] = 8'h72;
frames[12][3][0] = 8'h20;
frames[12][3][1] = 8'h44;
frames[12][3][2] = 8'h48;
frames[12][3][3] = 8'h68;
frames[12][3][4] = 8'h44;
frames[12][3][5] = 8'h44;
frames[12][3][6] = 8'h64;
frames[12][3][7] = 8'h68;
frames[12][3][8] = 8'h68;
frames[12][3][9] = 8'h89;
frames[12][3][10] = 8'had;
frames[12][3][11] = 8'had;
frames[12][3][12] = 8'had;
frames[12][3][13] = 8'had;
frames[12][3][14] = 8'had;
frames[12][3][15] = 8'had;
frames[12][3][16] = 8'had;
frames[12][3][17] = 8'h88;
frames[12][3][18] = 8'h89;
frames[12][3][19] = 8'h89;
frames[12][3][20] = 8'h64;
frames[12][3][21] = 8'h88;
frames[12][3][22] = 8'h89;
frames[12][3][23] = 8'had;
frames[12][3][24] = 8'h89;
frames[12][3][25] = 8'h64;
frames[12][3][26] = 8'ha9;
frames[12][3][27] = 8'had;
frames[12][3][28] = 8'h64;
frames[12][3][29] = 8'h64;
frames[12][3][30] = 8'h89;
frames[12][3][31] = 8'h88;
frames[12][3][32] = 8'h44;
frames[12][3][33] = 8'h24;
frames[12][3][34] = 8'h24;
frames[12][3][35] = 8'h44;
frames[12][3][36] = 8'h8d;
frames[12][3][37] = 8'h69;
frames[12][3][38] = 8'h4d;
frames[12][3][39] = 8'h92;
frames[12][4][0] = 8'h44;
frames[12][4][1] = 8'h48;
frames[12][4][2] = 8'h44;
frames[12][4][3] = 8'h44;
frames[12][4][4] = 8'h24;
frames[12][4][5] = 8'h00;
frames[12][4][6] = 8'h20;
frames[12][4][7] = 8'h24;
frames[12][4][8] = 8'h24;
frames[12][4][9] = 8'h44;
frames[12][4][10] = 8'h64;
frames[12][4][11] = 8'h89;
frames[12][4][12] = 8'had;
frames[12][4][13] = 8'had;
frames[12][4][14] = 8'had;
frames[12][4][15] = 8'had;
frames[12][4][16] = 8'had;
frames[12][4][17] = 8'h88;
frames[12][4][18] = 8'h88;
frames[12][4][19] = 8'h89;
frames[12][4][20] = 8'h88;
frames[12][4][21] = 8'h64;
frames[12][4][22] = 8'h89;
frames[12][4][23] = 8'h89;
frames[12][4][24] = 8'had;
frames[12][4][25] = 8'h88;
frames[12][4][26] = 8'h84;
frames[12][4][27] = 8'ha9;
frames[12][4][28] = 8'h89;
frames[12][4][29] = 8'h64;
frames[12][4][30] = 8'h44;
frames[12][4][31] = 8'h44;
frames[12][4][32] = 8'h44;
frames[12][4][33] = 8'h44;
frames[12][4][34] = 8'h44;
frames[12][4][35] = 8'h44;
frames[12][4][36] = 8'hb1;
frames[12][4][37] = 8'h8d;
frames[12][4][38] = 8'h91;
frames[12][4][39] = 8'h8d;
frames[12][5][0] = 8'h48;
frames[12][5][1] = 8'h44;
frames[12][5][2] = 8'h24;
frames[12][5][3] = 8'h24;
frames[12][5][4] = 8'h00;
frames[12][5][5] = 8'h00;
frames[12][5][6] = 8'h00;
frames[12][5][7] = 8'h24;
frames[12][5][8] = 8'h24;
frames[12][5][9] = 8'h20;
frames[12][5][10] = 8'h20;
frames[12][5][11] = 8'h44;
frames[12][5][12] = 8'had;
frames[12][5][13] = 8'had;
frames[12][5][14] = 8'had;
frames[12][5][15] = 8'had;
frames[12][5][16] = 8'had;
frames[12][5][17] = 8'h68;
frames[12][5][18] = 8'h64;
frames[12][5][19] = 8'h89;
frames[12][5][20] = 8'h89;
frames[12][5][21] = 8'h68;
frames[12][5][22] = 8'h88;
frames[12][5][23] = 8'h89;
frames[12][5][24] = 8'had;
frames[12][5][25] = 8'had;
frames[12][5][26] = 8'h84;
frames[12][5][27] = 8'ha9;
frames[12][5][28] = 8'had;
frames[12][5][29] = 8'h64;
frames[12][5][30] = 8'h44;
frames[12][5][31] = 8'h64;
frames[12][5][32] = 8'h64;
frames[12][5][33] = 8'h64;
frames[12][5][34] = 8'h64;
frames[12][5][35] = 8'h64;
frames[12][5][36] = 8'h68;
frames[12][5][37] = 8'hb1;
frames[12][5][38] = 8'hb1;
frames[12][5][39] = 8'h64;
frames[12][6][0] = 8'h24;
frames[12][6][1] = 8'h24;
frames[12][6][2] = 8'h44;
frames[12][6][3] = 8'h24;
frames[12][6][4] = 8'h24;
frames[12][6][5] = 8'h20;
frames[12][6][6] = 8'h44;
frames[12][6][7] = 8'h8d;
frames[12][6][8] = 8'h6d;
frames[12][6][9] = 8'h48;
frames[12][6][10] = 8'h24;
frames[12][6][11] = 8'h24;
frames[12][6][12] = 8'h44;
frames[12][6][13] = 8'h8d;
frames[12][6][14] = 8'had;
frames[12][6][15] = 8'had;
frames[12][6][16] = 8'h88;
frames[12][6][17] = 8'h64;
frames[12][6][18] = 8'h64;
frames[12][6][19] = 8'h88;
frames[12][6][20] = 8'h89;
frames[12][6][21] = 8'ha9;
frames[12][6][22] = 8'h64;
frames[12][6][23] = 8'h88;
frames[12][6][24] = 8'h88;
frames[12][6][25] = 8'had;
frames[12][6][26] = 8'h88;
frames[12][6][27] = 8'h88;
frames[12][6][28] = 8'had;
frames[12][6][29] = 8'h88;
frames[12][6][30] = 8'h64;
frames[12][6][31] = 8'h64;
frames[12][6][32] = 8'h64;
frames[12][6][33] = 8'h64;
frames[12][6][34] = 8'h64;
frames[12][6][35] = 8'h64;
frames[12][6][36] = 8'h64;
frames[12][6][37] = 8'h64;
frames[12][6][38] = 8'h64;
frames[12][6][39] = 8'h68;
frames[12][7][0] = 8'h6d;
frames[12][7][1] = 8'h6d;
frames[12][7][2] = 8'h8d;
frames[12][7][3] = 8'h8d;
frames[12][7][4] = 8'h8d;
frames[12][7][5] = 8'h8d;
frames[12][7][6] = 8'h8d;
frames[12][7][7] = 8'h91;
frames[12][7][8] = 8'h91;
frames[12][7][9] = 8'hb1;
frames[12][7][10] = 8'h8d;
frames[12][7][11] = 8'h68;
frames[12][7][12] = 8'h68;
frames[12][7][13] = 8'h68;
frames[12][7][14] = 8'h8d;
frames[12][7][15] = 8'h89;
frames[12][7][16] = 8'h88;
frames[12][7][17] = 8'h64;
frames[12][7][18] = 8'h64;
frames[12][7][19] = 8'h64;
frames[12][7][20] = 8'h88;
frames[12][7][21] = 8'ha9;
frames[12][7][22] = 8'h89;
frames[12][7][23] = 8'h64;
frames[12][7][24] = 8'h88;
frames[12][7][25] = 8'h89;
frames[12][7][26] = 8'had;
frames[12][7][27] = 8'h84;
frames[12][7][28] = 8'had;
frames[12][7][29] = 8'h89;
frames[12][7][30] = 8'h44;
frames[12][7][31] = 8'h44;
frames[12][7][32] = 8'h44;
frames[12][7][33] = 8'h44;
frames[12][7][34] = 8'h64;
frames[12][7][35] = 8'h68;
frames[12][7][36] = 8'h68;
frames[12][7][37] = 8'h68;
frames[12][7][38] = 8'h68;
frames[12][7][39] = 8'h68;
frames[12][8][0] = 8'hb1;
frames[12][8][1] = 8'hb1;
frames[12][8][2] = 8'hb1;
frames[12][8][3] = 8'hb1;
frames[12][8][4] = 8'hb1;
frames[12][8][5] = 8'hb1;
frames[12][8][6] = 8'hb1;
frames[12][8][7] = 8'hb1;
frames[12][8][8] = 8'hb1;
frames[12][8][9] = 8'hb1;
frames[12][8][10] = 8'h8d;
frames[12][8][11] = 8'h8d;
frames[12][8][12] = 8'h8d;
frames[12][8][13] = 8'h6c;
frames[12][8][14] = 8'h8d;
frames[12][8][15] = 8'h68;
frames[12][8][16] = 8'h64;
frames[12][8][17] = 8'h64;
frames[12][8][18] = 8'h64;
frames[12][8][19] = 8'h64;
frames[12][8][20] = 8'h64;
frames[12][8][21] = 8'h88;
frames[12][8][22] = 8'h89;
frames[12][8][23] = 8'h64;
frames[12][8][24] = 8'h64;
frames[12][8][25] = 8'h89;
frames[12][8][26] = 8'had;
frames[12][8][27] = 8'h84;
frames[12][8][28] = 8'h89;
frames[12][8][29] = 8'ha9;
frames[12][8][30] = 8'h24;
frames[12][8][31] = 8'h24;
frames[12][8][32] = 8'h24;
frames[12][8][33] = 8'h24;
frames[12][8][34] = 8'h44;
frames[12][8][35] = 8'h44;
frames[12][8][36] = 8'h44;
frames[12][8][37] = 8'h44;
frames[12][8][38] = 8'h44;
frames[12][8][39] = 8'h44;
frames[12][9][0] = 8'h8d;
frames[12][9][1] = 8'h8d;
frames[12][9][2] = 8'h88;
frames[12][9][3] = 8'h88;
frames[12][9][4] = 8'h8d;
frames[12][9][5] = 8'h8d;
frames[12][9][6] = 8'had;
frames[12][9][7] = 8'h88;
frames[12][9][8] = 8'h84;
frames[12][9][9] = 8'h64;
frames[12][9][10] = 8'h64;
frames[12][9][11] = 8'had;
frames[12][9][12] = 8'hb1;
frames[12][9][13] = 8'hb1;
frames[12][9][14] = 8'h8d;
frames[12][9][15] = 8'h8d;
frames[12][9][16] = 8'h48;
frames[12][9][17] = 8'h24;
frames[12][9][18] = 8'h44;
frames[12][9][19] = 8'h64;
frames[12][9][20] = 8'h64;
frames[12][9][21] = 8'h68;
frames[12][9][22] = 8'h68;
frames[12][9][23] = 8'h89;
frames[12][9][24] = 8'h64;
frames[12][9][25] = 8'h88;
frames[12][9][26] = 8'had;
frames[12][9][27] = 8'h88;
frames[12][9][28] = 8'h84;
frames[12][9][29] = 8'ha9;
frames[12][9][30] = 8'h44;
frames[12][9][31] = 8'h24;
frames[12][9][32] = 8'h24;
frames[12][9][33] = 8'h24;
frames[12][9][34] = 8'h24;
frames[12][9][35] = 8'h24;
frames[12][9][36] = 8'h24;
frames[12][9][37] = 8'h24;
frames[12][9][38] = 8'h24;
frames[12][9][39] = 8'h24;
frames[12][10][0] = 8'h8d;
frames[12][10][1] = 8'h88;
frames[12][10][2] = 8'h84;
frames[12][10][3] = 8'h88;
frames[12][10][4] = 8'hb1;
frames[12][10][5] = 8'hb1;
frames[12][10][6] = 8'ha8;
frames[12][10][7] = 8'h64;
frames[12][10][8] = 8'h84;
frames[12][10][9] = 8'h84;
frames[12][10][10] = 8'h68;
frames[12][10][11] = 8'hd1;
frames[12][10][12] = 8'hd6;
frames[12][10][13] = 8'hb1;
frames[12][10][14] = 8'h8d;
frames[12][10][15] = 8'h91;
frames[12][10][16] = 8'h8d;
frames[12][10][17] = 8'h44;
frames[12][10][18] = 8'h44;
frames[12][10][19] = 8'h44;
frames[12][10][20] = 8'h64;
frames[12][10][21] = 8'h64;
frames[12][10][22] = 8'h64;
frames[12][10][23] = 8'h88;
frames[12][10][24] = 8'h88;
frames[12][10][25] = 8'h64;
frames[12][10][26] = 8'ha9;
frames[12][10][27] = 8'ha9;
frames[12][10][28] = 8'h84;
frames[12][10][29] = 8'ha9;
frames[12][10][30] = 8'h68;
frames[12][10][31] = 8'h20;
frames[12][10][32] = 8'h24;
frames[12][10][33] = 8'h24;
frames[12][10][34] = 8'h24;
frames[12][10][35] = 8'h24;
frames[12][10][36] = 8'h24;
frames[12][10][37] = 8'h24;
frames[12][10][38] = 8'h24;
frames[12][10][39] = 8'h24;
frames[12][11][0] = 8'h88;
frames[12][11][1] = 8'h88;
frames[12][11][2] = 8'h84;
frames[12][11][3] = 8'h84;
frames[12][11][4] = 8'h88;
frames[12][11][5] = 8'hb1;
frames[12][11][6] = 8'had;
frames[12][11][7] = 8'h88;
frames[12][11][8] = 8'ha8;
frames[12][11][9] = 8'h84;
frames[12][11][10] = 8'h88;
frames[12][11][11] = 8'hd1;
frames[12][11][12] = 8'hb5;
frames[12][11][13] = 8'hd5;
frames[12][11][14] = 8'hd6;
frames[12][11][15] = 8'hb6;
frames[12][11][16] = 8'hb2;
frames[12][11][17] = 8'h44;
frames[12][11][18] = 8'h44;
frames[12][11][19] = 8'h44;
frames[12][11][20] = 8'h44;
frames[12][11][21] = 8'h64;
frames[12][11][22] = 8'h64;
frames[12][11][23] = 8'h88;
frames[12][11][24] = 8'h88;
frames[12][11][25] = 8'h64;
frames[12][11][26] = 8'h88;
frames[12][11][27] = 8'ha9;
frames[12][11][28] = 8'h84;
frames[12][11][29] = 8'ha9;
frames[12][11][30] = 8'h68;
frames[12][11][31] = 8'h20;
frames[12][11][32] = 8'h24;
frames[12][11][33] = 8'h24;
frames[12][11][34] = 8'h24;
frames[12][11][35] = 8'h24;
frames[12][11][36] = 8'h24;
frames[12][11][37] = 8'h24;
frames[12][11][38] = 8'h24;
frames[12][11][39] = 8'h24;
frames[12][12][0] = 8'hcd;
frames[12][12][1] = 8'h84;
frames[12][12][2] = 8'ha4;
frames[12][12][3] = 8'h80;
frames[12][12][4] = 8'h88;
frames[12][12][5] = 8'hcd;
frames[12][12][6] = 8'hb1;
frames[12][12][7] = 8'hb1;
frames[12][12][8] = 8'had;
frames[12][12][9] = 8'h88;
frames[12][12][10] = 8'h84;
frames[12][12][11] = 8'ha8;
frames[12][12][12] = 8'h88;
frames[12][12][13] = 8'hd1;
frames[12][12][14] = 8'hd6;
frames[12][12][15] = 8'hd6;
frames[12][12][16] = 8'h91;
frames[12][12][17] = 8'h44;
frames[12][12][18] = 8'h44;
frames[12][12][19] = 8'h44;
frames[12][12][20] = 8'h44;
frames[12][12][21] = 8'h44;
frames[12][12][22] = 8'h44;
frames[12][12][23] = 8'h44;
frames[12][12][24] = 8'h64;
frames[12][12][25] = 8'h64;
frames[12][12][26] = 8'h84;
frames[12][12][27] = 8'h88;
frames[12][12][28] = 8'h84;
frames[12][12][29] = 8'h84;
frames[12][12][30] = 8'h44;
frames[12][12][31] = 8'h24;
frames[12][12][32] = 8'h24;
frames[12][12][33] = 8'h24;
frames[12][12][34] = 8'h24;
frames[12][12][35] = 8'h24;
frames[12][12][36] = 8'h24;
frames[12][12][37] = 8'h24;
frames[12][12][38] = 8'h24;
frames[12][12][39] = 8'h24;
frames[12][13][0] = 8'hf6;
frames[12][13][1] = 8'hac;
frames[12][13][2] = 8'ha4;
frames[12][13][3] = 8'h84;
frames[12][13][4] = 8'h84;
frames[12][13][5] = 8'ha8;
frames[12][13][6] = 8'h88;
frames[12][13][7] = 8'had;
frames[12][13][8] = 8'hd5;
frames[12][13][9] = 8'hb1;
frames[12][13][10] = 8'hd1;
frames[12][13][11] = 8'had;
frames[12][13][12] = 8'h88;
frames[12][13][13] = 8'hd1;
frames[12][13][14] = 8'hb1;
frames[12][13][15] = 8'hb6;
frames[12][13][16] = 8'h69;
frames[12][13][17] = 8'h44;
frames[12][13][18] = 8'h44;
frames[12][13][19] = 8'h44;
frames[12][13][20] = 8'h44;
frames[12][13][21] = 8'h44;
frames[12][13][22] = 8'h44;
frames[12][13][23] = 8'h44;
frames[12][13][24] = 8'h44;
frames[12][13][25] = 8'h48;
frames[12][13][26] = 8'h64;
frames[12][13][27] = 8'h88;
frames[12][13][28] = 8'h89;
frames[12][13][29] = 8'h64;
frames[12][13][30] = 8'h24;
frames[12][13][31] = 8'h24;
frames[12][13][32] = 8'h24;
frames[12][13][33] = 8'h24;
frames[12][13][34] = 8'h24;
frames[12][13][35] = 8'h24;
frames[12][13][36] = 8'h24;
frames[12][13][37] = 8'h24;
frames[12][13][38] = 8'h24;
frames[12][13][39] = 8'h24;
frames[12][14][0] = 8'hb1;
frames[12][14][1] = 8'hd5;
frames[12][14][2] = 8'ha8;
frames[12][14][3] = 8'h64;
frames[12][14][4] = 8'h84;
frames[12][14][5] = 8'h84;
frames[12][14][6] = 8'h88;
frames[12][14][7] = 8'had;
frames[12][14][8] = 8'hb1;
frames[12][14][9] = 8'hb1;
frames[12][14][10] = 8'hd6;
frames[12][14][11] = 8'hda;
frames[12][14][12] = 8'hb1;
frames[12][14][13] = 8'hb1;
frames[12][14][14] = 8'hb2;
frames[12][14][15] = 8'h6d;
frames[12][14][16] = 8'h44;
frames[12][14][17] = 8'h44;
frames[12][14][18] = 8'h44;
frames[12][14][19] = 8'h44;
frames[12][14][20] = 8'h48;
frames[12][14][21] = 8'h44;
frames[12][14][22] = 8'h48;
frames[12][14][23] = 8'h69;
frames[12][14][24] = 8'h8d;
frames[12][14][25] = 8'h69;
frames[12][14][26] = 8'h64;
frames[12][14][27] = 8'h89;
frames[12][14][28] = 8'had;
frames[12][14][29] = 8'h88;
frames[12][14][30] = 8'h88;
frames[12][14][31] = 8'h88;
frames[12][14][32] = 8'h48;
frames[12][14][33] = 8'h48;
frames[12][14][34] = 8'h48;
frames[12][14][35] = 8'h44;
frames[12][14][36] = 8'h24;
frames[12][14][37] = 8'h24;
frames[12][14][38] = 8'h24;
frames[12][14][39] = 8'h24;
frames[12][15][0] = 8'h88;
frames[12][15][1] = 8'hb1;
frames[12][15][2] = 8'hd1;
frames[12][15][3] = 8'hac;
frames[12][15][4] = 8'h88;
frames[12][15][5] = 8'h88;
frames[12][15][6] = 8'h8c;
frames[12][15][7] = 8'hb1;
frames[12][15][8] = 8'hb1;
frames[12][15][9] = 8'hb1;
frames[12][15][10] = 8'hd5;
frames[12][15][11] = 8'hd5;
frames[12][15][12] = 8'hb1;
frames[12][15][13] = 8'h91;
frames[12][15][14] = 8'h69;
frames[12][15][15] = 8'h24;
frames[12][15][16] = 8'h24;
frames[12][15][17] = 8'h44;
frames[12][15][18] = 8'h44;
frames[12][15][19] = 8'h6d;
frames[12][15][20] = 8'hb1;
frames[12][15][21] = 8'h88;
frames[12][15][22] = 8'h88;
frames[12][15][23] = 8'h8d;
frames[12][15][24] = 8'had;
frames[12][15][25] = 8'had;
frames[12][15][26] = 8'had;
frames[12][15][27] = 8'hb1;
frames[12][15][28] = 8'hd1;
frames[12][15][29] = 8'hd1;
frames[12][15][30] = 8'hb1;
frames[12][15][31] = 8'hb1;
frames[12][15][32] = 8'hb1;
frames[12][15][33] = 8'hb1;
frames[12][15][34] = 8'hb1;
frames[12][15][35] = 8'h68;
frames[12][15][36] = 8'h48;
frames[12][15][37] = 8'h6d;
frames[12][15][38] = 8'h24;
frames[12][15][39] = 8'h24;
frames[12][16][0] = 8'h8d;
frames[12][16][1] = 8'hd6;
frames[12][16][2] = 8'hd6;
frames[12][16][3] = 8'hd5;
frames[12][16][4] = 8'hb1;
frames[12][16][5] = 8'h8d;
frames[12][16][6] = 8'had;
frames[12][16][7] = 8'hd1;
frames[12][16][8] = 8'hb1;
frames[12][16][9] = 8'hb1;
frames[12][16][10] = 8'hb1;
frames[12][16][11] = 8'hb1;
frames[12][16][12] = 8'h68;
frames[12][16][13] = 8'h44;
frames[12][16][14] = 8'h24;
frames[12][16][15] = 8'h44;
frames[12][16][16] = 8'h48;
frames[12][16][17] = 8'h69;
frames[12][16][18] = 8'had;
frames[12][16][19] = 8'had;
frames[12][16][20] = 8'hb1;
frames[12][16][21] = 8'hd1;
frames[12][16][22] = 8'h8c;
frames[12][16][23] = 8'h8c;
frames[12][16][24] = 8'h88;
frames[12][16][25] = 8'hb1;
frames[12][16][26] = 8'hd1;
frames[12][16][27] = 8'hd5;
frames[12][16][28] = 8'hd5;
frames[12][16][29] = 8'hd1;
frames[12][16][30] = 8'had;
frames[12][16][31] = 8'h88;
frames[12][16][32] = 8'h88;
frames[12][16][33] = 8'ha8;
frames[12][16][34] = 8'had;
frames[12][16][35] = 8'hd1;
frames[12][16][36] = 8'hb1;
frames[12][16][37] = 8'hb1;
frames[12][16][38] = 8'h48;
frames[12][16][39] = 8'h44;
frames[12][17][0] = 8'hd6;
frames[12][17][1] = 8'hd6;
frames[12][17][2] = 8'hb5;
frames[12][17][3] = 8'hb1;
frames[12][17][4] = 8'hd6;
frames[12][17][5] = 8'hb1;
frames[12][17][6] = 8'hb1;
frames[12][17][7] = 8'hd5;
frames[12][17][8] = 8'hb6;
frames[12][17][9] = 8'h91;
frames[12][17][10] = 8'h48;
frames[12][17][11] = 8'h20;
frames[12][17][12] = 8'h20;
frames[12][17][13] = 8'h20;
frames[12][17][14] = 8'h48;
frames[12][17][15] = 8'h8d;
frames[12][17][16] = 8'h88;
frames[12][17][17] = 8'h88;
frames[12][17][18] = 8'h88;
frames[12][17][19] = 8'ha8;
frames[12][17][20] = 8'hb1;
frames[12][17][21] = 8'hb1;
frames[12][17][22] = 8'h8d;
frames[12][17][23] = 8'hb1;
frames[12][17][24] = 8'hd1;
frames[12][17][25] = 8'hd5;
frames[12][17][26] = 8'hd5;
frames[12][17][27] = 8'hd5;
frames[12][17][28] = 8'hd5;
frames[12][17][29] = 8'hb1;
frames[12][17][30] = 8'hd6;
frames[12][17][31] = 8'hd1;
frames[12][17][32] = 8'hb1;
frames[12][17][33] = 8'hb1;
frames[12][17][34] = 8'hb1;
frames[12][17][35] = 8'hd1;
frames[12][17][36] = 8'hb5;
frames[12][17][37] = 8'hb5;
frames[12][17][38] = 8'h91;
frames[12][17][39] = 8'h6d;
frames[12][18][0] = 8'hda;
frames[12][18][1] = 8'hd6;
frames[12][18][2] = 8'hb5;
frames[12][18][3] = 8'hd6;
frames[12][18][4] = 8'hd6;
frames[12][18][5] = 8'hb1;
frames[12][18][6] = 8'h91;
frames[12][18][7] = 8'h6d;
frames[12][18][8] = 8'h44;
frames[12][18][9] = 8'h20;
frames[12][18][10] = 8'h20;
frames[12][18][11] = 8'h20;
frames[12][18][12] = 8'h20;
frames[12][18][13] = 8'h48;
frames[12][18][14] = 8'hb1;
frames[12][18][15] = 8'hb1;
frames[12][18][16] = 8'had;
frames[12][18][17] = 8'ha8;
frames[12][18][18] = 8'ha4;
frames[12][18][19] = 8'ha4;
frames[12][18][20] = 8'hd1;
frames[12][18][21] = 8'hb1;
frames[12][18][22] = 8'had;
frames[12][18][23] = 8'hb1;
frames[12][18][24] = 8'hd5;
frames[12][18][25] = 8'hd5;
frames[12][18][26] = 8'hd6;
frames[12][18][27] = 8'hd5;
frames[12][18][28] = 8'hda;
frames[12][18][29] = 8'hd5;
frames[12][18][30] = 8'hd1;
frames[12][18][31] = 8'hd5;
frames[12][18][32] = 8'hb1;
frames[12][18][33] = 8'hd5;
frames[12][18][34] = 8'hd6;
frames[12][18][35] = 8'hd6;
frames[12][18][36] = 8'hd6;
frames[12][18][37] = 8'hb1;
frames[12][18][38] = 8'h91;
frames[12][18][39] = 8'h91;
frames[12][19][0] = 8'h8d;
frames[12][19][1] = 8'h8d;
frames[12][19][2] = 8'h8d;
frames[12][19][3] = 8'h6d;
frames[12][19][4] = 8'h48;
frames[12][19][5] = 8'h44;
frames[12][19][6] = 8'h24;
frames[12][19][7] = 8'h24;
frames[12][19][8] = 8'h24;
frames[12][19][9] = 8'h24;
frames[12][19][10] = 8'h24;
frames[12][19][11] = 8'h24;
frames[12][19][12] = 8'h69;
frames[12][19][13] = 8'hb1;
frames[12][19][14] = 8'hd6;
frames[12][19][15] = 8'hd6;
frames[12][19][16] = 8'hcd;
frames[12][19][17] = 8'h88;
frames[12][19][18] = 8'h84;
frames[12][19][19] = 8'ha4;
frames[12][19][20] = 8'hb1;
frames[12][19][21] = 8'hd1;
frames[12][19][22] = 8'had;
frames[12][19][23] = 8'had;
frames[12][19][24] = 8'hd5;
frames[12][19][25] = 8'hd6;
frames[12][19][26] = 8'hd6;
frames[12][19][27] = 8'hb1;
frames[12][19][28] = 8'hd6;
frames[12][19][29] = 8'hd5;
frames[12][19][30] = 8'ha8;
frames[12][19][31] = 8'h88;
frames[12][19][32] = 8'h88;
frames[12][19][33] = 8'ha8;
frames[12][19][34] = 8'had;
frames[12][19][35] = 8'hd6;
frames[12][19][36] = 8'hd6;
frames[12][19][37] = 8'hb1;
frames[12][19][38] = 8'hb1;
frames[12][19][39] = 8'h91;
frames[12][20][0] = 8'h24;
frames[12][20][1] = 8'h24;
frames[12][20][2] = 8'h24;
frames[12][20][3] = 8'h24;
frames[12][20][4] = 8'h24;
frames[12][20][5] = 8'h24;
frames[12][20][6] = 8'h24;
frames[12][20][7] = 8'h24;
frames[12][20][8] = 8'h24;
frames[12][20][9] = 8'h24;
frames[12][20][10] = 8'h24;
frames[12][20][11] = 8'h44;
frames[12][20][12] = 8'h91;
frames[12][20][13] = 8'hb1;
frames[12][20][14] = 8'hd6;
frames[12][20][15] = 8'hd1;
frames[12][20][16] = 8'ha4;
frames[12][20][17] = 8'ha4;
frames[12][20][18] = 8'ha4;
frames[12][20][19] = 8'ha4;
frames[12][20][20] = 8'had;
frames[12][20][21] = 8'hb1;
frames[12][20][22] = 8'hcd;
frames[12][20][23] = 8'ha8;
frames[12][20][24] = 8'ha8;
frames[12][20][25] = 8'hcd;
frames[12][20][26] = 8'hd1;
frames[12][20][27] = 8'hb1;
frames[12][20][28] = 8'hd5;
frames[12][20][29] = 8'had;
frames[12][20][30] = 8'h84;
frames[12][20][31] = 8'ha4;
frames[12][20][32] = 8'ha4;
frames[12][20][33] = 8'ha4;
frames[12][20][34] = 8'h88;
frames[12][20][35] = 8'hd1;
frames[12][20][36] = 8'hd6;
frames[12][20][37] = 8'hd6;
frames[12][20][38] = 8'hb1;
frames[12][20][39] = 8'hb1;
frames[12][21][0] = 8'h48;
frames[12][21][1] = 8'h44;
frames[12][21][2] = 8'h24;
frames[12][21][3] = 8'h24;
frames[12][21][4] = 8'h24;
frames[12][21][5] = 8'h44;
frames[12][21][6] = 8'h24;
frames[12][21][7] = 8'h24;
frames[12][21][8] = 8'h24;
frames[12][21][9] = 8'h24;
frames[12][21][10] = 8'h24;
frames[12][21][11] = 8'h24;
frames[12][21][12] = 8'h91;
frames[12][21][13] = 8'h91;
frames[12][21][14] = 8'hd1;
frames[12][21][15] = 8'hb1;
frames[12][21][16] = 8'ha8;
frames[12][21][17] = 8'ha8;
frames[12][21][18] = 8'hcd;
frames[12][21][19] = 8'hd1;
frames[12][21][20] = 8'hb1;
frames[12][21][21] = 8'h8d;
frames[12][21][22] = 8'hd1;
frames[12][21][23] = 8'hd1;
frames[12][21][24] = 8'hc8;
frames[12][21][25] = 8'ha8;
frames[12][21][26] = 8'ha8;
frames[12][21][27] = 8'ha8;
frames[12][21][28] = 8'hb1;
frames[12][21][29] = 8'hb1;
frames[12][21][30] = 8'ha4;
frames[12][21][31] = 8'h84;
frames[12][21][32] = 8'h84;
frames[12][21][33] = 8'ha4;
frames[12][21][34] = 8'had;
frames[12][21][35] = 8'hd1;
frames[12][21][36] = 8'hb1;
frames[12][21][37] = 8'hb1;
frames[12][21][38] = 8'h8d;
frames[12][21][39] = 8'h68;
frames[12][22][0] = 8'h49;
frames[12][22][1] = 8'h48;
frames[12][22][2] = 8'h48;
frames[12][22][3] = 8'h44;
frames[12][22][4] = 8'h24;
frames[12][22][5] = 8'h24;
frames[12][22][6] = 8'h24;
frames[12][22][7] = 8'h24;
frames[12][22][8] = 8'h24;
frames[12][22][9] = 8'h24;
frames[12][22][10] = 8'h24;
frames[12][22][11] = 8'h24;
frames[12][22][12] = 8'h69;
frames[12][22][13] = 8'hb1;
frames[12][22][14] = 8'hb1;
frames[12][22][15] = 8'hd1;
frames[12][22][16] = 8'hd5;
frames[12][22][17] = 8'hd1;
frames[12][22][18] = 8'had;
frames[12][22][19] = 8'hd5;
frames[12][22][20] = 8'hb5;
frames[12][22][21] = 8'hb1;
frames[12][22][22] = 8'hd5;
frames[12][22][23] = 8'hb1;
frames[12][22][24] = 8'hd1;
frames[12][22][25] = 8'hac;
frames[12][22][26] = 8'ha8;
frames[12][22][27] = 8'had;
frames[12][22][28] = 8'hb1;
frames[12][22][29] = 8'hb1;
frames[12][22][30] = 8'had;
frames[12][22][31] = 8'hac;
frames[12][22][32] = 8'hac;
frames[12][22][33] = 8'hd1;
frames[12][22][34] = 8'hd6;
frames[12][22][35] = 8'hb1;
frames[12][22][36] = 8'hb6;
frames[12][22][37] = 8'h8d;
frames[12][22][38] = 8'h24;
frames[12][22][39] = 8'h24;
frames[12][23][0] = 8'h44;
frames[12][23][1] = 8'h48;
frames[12][23][2] = 8'h48;
frames[12][23][3] = 8'h69;
frames[12][23][4] = 8'h49;
frames[12][23][5] = 8'h48;
frames[12][23][6] = 8'h44;
frames[12][23][7] = 8'h24;
frames[12][23][8] = 8'h24;
frames[12][23][9] = 8'h24;
frames[12][23][10] = 8'h24;
frames[12][23][11] = 8'h24;
frames[12][23][12] = 8'h24;
frames[12][23][13] = 8'h6d;
frames[12][23][14] = 8'hb1;
frames[12][23][15] = 8'hb2;
frames[12][23][16] = 8'hd6;
frames[12][23][17] = 8'hd6;
frames[12][23][18] = 8'hd6;
frames[12][23][19] = 8'hd6;
frames[12][23][20] = 8'hd5;
frames[12][23][21] = 8'hd5;
frames[12][23][22] = 8'hd6;
frames[12][23][23] = 8'hd5;
frames[12][23][24] = 8'hd6;
frames[12][23][25] = 8'hd6;
frames[12][23][26] = 8'hd6;
frames[12][23][27] = 8'hd6;
frames[12][23][28] = 8'hd5;
frames[12][23][29] = 8'hd5;
frames[12][23][30] = 8'hfa;
frames[12][23][31] = 8'hd6;
frames[12][23][32] = 8'hd5;
frames[12][23][33] = 8'hb1;
frames[12][23][34] = 8'hb1;
frames[12][23][35] = 8'h6c;
frames[12][23][36] = 8'h44;
frames[12][23][37] = 8'h24;
frames[12][23][38] = 8'h44;
frames[12][23][39] = 8'h48;
frames[12][24][0] = 8'h68;
frames[12][24][1] = 8'h48;
frames[12][24][2] = 8'h44;
frames[12][24][3] = 8'h44;
frames[12][24][4] = 8'h44;
frames[12][24][5] = 8'h44;
frames[12][24][6] = 8'h49;
frames[12][24][7] = 8'h49;
frames[12][24][8] = 8'h48;
frames[12][24][9] = 8'h44;
frames[12][24][10] = 8'h24;
frames[12][24][11] = 8'h24;
frames[12][24][12] = 8'h24;
frames[12][24][13] = 8'h24;
frames[12][24][14] = 8'h44;
frames[12][24][15] = 8'h6d;
frames[12][24][16] = 8'hb1;
frames[12][24][17] = 8'hd6;
frames[12][24][18] = 8'hd6;
frames[12][24][19] = 8'hd6;
frames[12][24][20] = 8'hd6;
frames[12][24][21] = 8'hd5;
frames[12][24][22] = 8'hd5;
frames[12][24][23] = 8'hd6;
frames[12][24][24] = 8'hd6;
frames[12][24][25] = 8'hd6;
frames[12][24][26] = 8'hd6;
frames[12][24][27] = 8'hd6;
frames[12][24][28] = 8'hd6;
frames[12][24][29] = 8'hb6;
frames[12][24][30] = 8'hb1;
frames[12][24][31] = 8'h8d;
frames[12][24][32] = 8'h69;
frames[12][24][33] = 8'h44;
frames[12][24][34] = 8'h24;
frames[12][24][35] = 8'h20;
frames[12][24][36] = 8'h24;
frames[12][24][37] = 8'h44;
frames[12][24][38] = 8'h48;
frames[12][24][39] = 8'h49;
frames[12][25][0] = 8'h8d;
frames[12][25][1] = 8'h8d;
frames[12][25][2] = 8'h8d;
frames[12][25][3] = 8'h68;
frames[12][25][4] = 8'h68;
frames[12][25][5] = 8'h44;
frames[12][25][6] = 8'h44;
frames[12][25][7] = 8'h44;
frames[12][25][8] = 8'h44;
frames[12][25][9] = 8'h44;
frames[12][25][10] = 8'h48;
frames[12][25][11] = 8'h48;
frames[12][25][12] = 8'h48;
frames[12][25][13] = 8'h44;
frames[12][25][14] = 8'h24;
frames[12][25][15] = 8'h24;
frames[12][25][16] = 8'h24;
frames[12][25][17] = 8'h24;
frames[12][25][18] = 8'h48;
frames[12][25][19] = 8'h48;
frames[12][25][20] = 8'h68;
frames[12][25][21] = 8'h68;
frames[12][25][22] = 8'h68;
frames[12][25][23] = 8'h68;
frames[12][25][24] = 8'h68;
frames[12][25][25] = 8'h48;
frames[12][25][26] = 8'h48;
frames[12][25][27] = 8'h44;
frames[12][25][28] = 8'h44;
frames[12][25][29] = 8'h44;
frames[12][25][30] = 8'h24;
frames[12][25][31] = 8'h20;
frames[12][25][32] = 8'h00;
frames[12][25][33] = 8'h00;
frames[12][25][34] = 8'h24;
frames[12][25][35] = 8'h44;
frames[12][25][36] = 8'h49;
frames[12][25][37] = 8'h49;
frames[12][25][38] = 8'h48;
frames[12][25][39] = 8'h48;
frames[12][26][0] = 8'hb1;
frames[12][26][1] = 8'hb1;
frames[12][26][2] = 8'hb1;
frames[12][26][3] = 8'had;
frames[12][26][4] = 8'h8c;
frames[12][26][5] = 8'h8c;
frames[12][26][6] = 8'h68;
frames[12][26][7] = 8'h64;
frames[12][26][8] = 8'h44;
frames[12][26][9] = 8'h44;
frames[12][26][10] = 8'h44;
frames[12][26][11] = 8'h44;
frames[12][26][12] = 8'h44;
frames[12][26][13] = 8'h48;
frames[12][26][14] = 8'h48;
frames[12][26][15] = 8'h48;
frames[12][26][16] = 8'h44;
frames[12][26][17] = 8'h24;
frames[12][26][18] = 8'h20;
frames[12][26][19] = 8'h00;
frames[12][26][20] = 8'h00;
frames[12][26][21] = 8'h00;
frames[12][26][22] = 8'h00;
frames[12][26][23] = 8'h00;
frames[12][26][24] = 8'h00;
frames[12][26][25] = 8'h00;
frames[12][26][26] = 8'h00;
frames[12][26][27] = 8'h00;
frames[12][26][28] = 8'h00;
frames[12][26][29] = 8'h00;
frames[12][26][30] = 8'h00;
frames[12][26][31] = 8'h00;
frames[12][26][32] = 8'h20;
frames[12][26][33] = 8'h24;
frames[12][26][34] = 8'h44;
frames[12][26][35] = 8'h49;
frames[12][26][36] = 8'h69;
frames[12][26][37] = 8'h48;
frames[12][26][38] = 8'h44;
frames[12][26][39] = 8'h44;
frames[12][27][0] = 8'hb1;
frames[12][27][1] = 8'hb1;
frames[12][27][2] = 8'hb1;
frames[12][27][3] = 8'hb1;
frames[12][27][4] = 8'hb1;
frames[12][27][5] = 8'had;
frames[12][27][6] = 8'had;
frames[12][27][7] = 8'h8c;
frames[12][27][8] = 8'h88;
frames[12][27][9] = 8'h68;
frames[12][27][10] = 8'h48;
frames[12][27][11] = 8'h44;
frames[12][27][12] = 8'h44;
frames[12][27][13] = 8'h44;
frames[12][27][14] = 8'h44;
frames[12][27][15] = 8'h44;
frames[12][27][16] = 8'h48;
frames[12][27][17] = 8'h48;
frames[12][27][18] = 8'h48;
frames[12][27][19] = 8'h44;
frames[12][27][20] = 8'h44;
frames[12][27][21] = 8'h24;
frames[12][27][22] = 8'h24;
frames[12][27][23] = 8'h24;
frames[12][27][24] = 8'h24;
frames[12][27][25] = 8'h24;
frames[12][27][26] = 8'h24;
frames[12][27][27] = 8'h24;
frames[12][27][28] = 8'h24;
frames[12][27][29] = 8'h24;
frames[12][27][30] = 8'h24;
frames[12][27][31] = 8'h24;
frames[12][27][32] = 8'h44;
frames[12][27][33] = 8'h49;
frames[12][27][34] = 8'h69;
frames[12][27][35] = 8'h69;
frames[12][27][36] = 8'h44;
frames[12][27][37] = 8'h44;
frames[12][27][38] = 8'h44;
frames[12][27][39] = 8'h44;
frames[12][28][0] = 8'hb1;
frames[12][28][1] = 8'hb1;
frames[12][28][2] = 8'hb1;
frames[12][28][3] = 8'hb1;
frames[12][28][4] = 8'hb1;
frames[12][28][5] = 8'hb1;
frames[12][28][6] = 8'hb1;
frames[12][28][7] = 8'had;
frames[12][28][8] = 8'had;
frames[12][28][9] = 8'hac;
frames[12][28][10] = 8'h8c;
frames[12][28][11] = 8'h8c;
frames[12][28][12] = 8'h68;
frames[12][28][13] = 8'h68;
frames[12][28][14] = 8'h44;
frames[12][28][15] = 8'h44;
frames[12][28][16] = 8'h44;
frames[12][28][17] = 8'h44;
frames[12][28][18] = 8'h44;
frames[12][28][19] = 8'h44;
frames[12][28][20] = 8'h48;
frames[12][28][21] = 8'h48;
frames[12][28][22] = 8'h44;
frames[12][28][23] = 8'h44;
frames[12][28][24] = 8'h44;
frames[12][28][25] = 8'h44;
frames[12][28][26] = 8'h24;
frames[12][28][27] = 8'h24;
frames[12][28][28] = 8'h24;
frames[12][28][29] = 8'h24;
frames[12][28][30] = 8'h44;
frames[12][28][31] = 8'h48;
frames[12][28][32] = 8'h69;
frames[12][28][33] = 8'h69;
frames[12][28][34] = 8'h44;
frames[12][28][35] = 8'h44;
frames[12][28][36] = 8'h44;
frames[12][28][37] = 8'h44;
frames[12][28][38] = 8'h44;
frames[12][28][39] = 8'h44;
frames[12][29][0] = 8'hb1;
frames[12][29][1] = 8'hb1;
frames[12][29][2] = 8'hb1;
frames[12][29][3] = 8'hb1;
frames[12][29][4] = 8'hb1;
frames[12][29][5] = 8'hb1;
frames[12][29][6] = 8'hb1;
frames[12][29][7] = 8'had;
frames[12][29][8] = 8'had;
frames[12][29][9] = 8'had;
frames[12][29][10] = 8'had;
frames[12][29][11] = 8'had;
frames[12][29][12] = 8'h8d;
frames[12][29][13] = 8'h8c;
frames[12][29][14] = 8'h88;
frames[12][29][15] = 8'h68;
frames[12][29][16] = 8'h48;
frames[12][29][17] = 8'h44;
frames[12][29][18] = 8'h44;
frames[12][29][19] = 8'h44;
frames[12][29][20] = 8'h44;
frames[12][29][21] = 8'h44;
frames[12][29][22] = 8'h44;
frames[12][29][23] = 8'h48;
frames[12][29][24] = 8'h48;
frames[12][29][25] = 8'h44;
frames[12][29][26] = 8'h44;
frames[12][29][27] = 8'h44;
frames[12][29][28] = 8'h44;
frames[12][29][29] = 8'h48;
frames[12][29][30] = 8'h69;
frames[12][29][31] = 8'h48;
frames[12][29][32] = 8'h44;
frames[12][29][33] = 8'h44;
frames[12][29][34] = 8'h44;
frames[12][29][35] = 8'h44;
frames[12][29][36] = 8'h44;
frames[12][29][37] = 8'h44;
frames[12][29][38] = 8'h44;
frames[12][29][39] = 8'h44;
frames[13][0][0] = 8'hd6;
frames[13][0][1] = 8'hfa;
frames[13][0][2] = 8'hfa;
frames[13][0][3] = 8'hfa;
frames[13][0][4] = 8'hfa;
frames[13][0][5] = 8'hfa;
frames[13][0][6] = 8'hfa;
frames[13][0][7] = 8'hb1;
frames[13][0][8] = 8'had;
frames[13][0][9] = 8'had;
frames[13][0][10] = 8'had;
frames[13][0][11] = 8'h88;
frames[13][0][12] = 8'had;
frames[13][0][13] = 8'h68;
frames[13][0][14] = 8'h40;
frames[13][0][15] = 8'h40;
frames[13][0][16] = 8'h68;
frames[13][0][17] = 8'hd6;
frames[13][0][18] = 8'hd5;
frames[13][0][19] = 8'hd5;
frames[13][0][20] = 8'hd5;
frames[13][0][21] = 8'hd5;
frames[13][0][22] = 8'hd5;
frames[13][0][23] = 8'hd5;
frames[13][0][24] = 8'hd5;
frames[13][0][25] = 8'hd5;
frames[13][0][26] = 8'hd5;
frames[13][0][27] = 8'hb1;
frames[13][0][28] = 8'h91;
frames[13][0][29] = 8'h69;
frames[13][0][30] = 8'h44;
frames[13][0][31] = 8'h24;
frames[13][0][32] = 8'h49;
frames[13][0][33] = 8'h6d;
frames[13][0][34] = 8'h8d;
frames[13][0][35] = 8'h8d;
frames[13][0][36] = 8'h69;
frames[13][0][37] = 8'h8d;
frames[13][0][38] = 8'h6d;
frames[13][0][39] = 8'h44;
frames[13][1][0] = 8'hda;
frames[13][1][1] = 8'hfa;
frames[13][1][2] = 8'hfa;
frames[13][1][3] = 8'hfa;
frames[13][1][4] = 8'hfa;
frames[13][1][5] = 8'hfa;
frames[13][1][6] = 8'hfa;
frames[13][1][7] = 8'hb1;
frames[13][1][8] = 8'had;
frames[13][1][9] = 8'had;
frames[13][1][10] = 8'had;
frames[13][1][11] = 8'h88;
frames[13][1][12] = 8'had;
frames[13][1][13] = 8'h68;
frames[13][1][14] = 8'h40;
frames[13][1][15] = 8'h44;
frames[13][1][16] = 8'had;
frames[13][1][17] = 8'hd6;
frames[13][1][18] = 8'hd5;
frames[13][1][19] = 8'hd5;
frames[13][1][20] = 8'hd6;
frames[13][1][21] = 8'hd6;
frames[13][1][22] = 8'hd5;
frames[13][1][23] = 8'hd5;
frames[13][1][24] = 8'hd5;
frames[13][1][25] = 8'hb1;
frames[13][1][26] = 8'h8d;
frames[13][1][27] = 8'h44;
frames[13][1][28] = 8'h24;
frames[13][1][29] = 8'h20;
frames[13][1][30] = 8'h20;
frames[13][1][31] = 8'h24;
frames[13][1][32] = 8'h20;
frames[13][1][33] = 8'h20;
frames[13][1][34] = 8'h24;
frames[13][1][35] = 8'h44;
frames[13][1][36] = 8'h92;
frames[13][1][37] = 8'hda;
frames[13][1][38] = 8'hda;
frames[13][1][39] = 8'h6d;
frames[13][2][0] = 8'hfa;
frames[13][2][1] = 8'hfa;
frames[13][2][2] = 8'hfa;
frames[13][2][3] = 8'hfa;
frames[13][2][4] = 8'hfa;
frames[13][2][5] = 8'hfa;
frames[13][2][6] = 8'hfa;
frames[13][2][7] = 8'hb1;
frames[13][2][8] = 8'had;
frames[13][2][9] = 8'had;
frames[13][2][10] = 8'had;
frames[13][2][11] = 8'h88;
frames[13][2][12] = 8'h8d;
frames[13][2][13] = 8'h88;
frames[13][2][14] = 8'h44;
frames[13][2][15] = 8'h64;
frames[13][2][16] = 8'hb1;
frames[13][2][17] = 8'hd5;
frames[13][2][18] = 8'hd5;
frames[13][2][19] = 8'hd5;
frames[13][2][20] = 8'hd5;
frames[13][2][21] = 8'hd6;
frames[13][2][22] = 8'hb6;
frames[13][2][23] = 8'hb1;
frames[13][2][24] = 8'h48;
frames[13][2][25] = 8'h24;
frames[13][2][26] = 8'h24;
frames[13][2][27] = 8'h20;
frames[13][2][28] = 8'h20;
frames[13][2][29] = 8'h00;
frames[13][2][30] = 8'h00;
frames[13][2][31] = 8'h20;
frames[13][2][32] = 8'h20;
frames[13][2][33] = 8'h20;
frames[13][2][34] = 8'h20;
frames[13][2][35] = 8'h20;
frames[13][2][36] = 8'h6e;
frames[13][2][37] = 8'h49;
frames[13][2][38] = 8'h4e;
frames[13][2][39] = 8'h92;
frames[13][3][0] = 8'hfa;
frames[13][3][1] = 8'hfa;
frames[13][3][2] = 8'hfa;
frames[13][3][3] = 8'hfa;
frames[13][3][4] = 8'hfa;
frames[13][3][5] = 8'hfa;
frames[13][3][6] = 8'hfa;
frames[13][3][7] = 8'had;
frames[13][3][8] = 8'had;
frames[13][3][9] = 8'had;
frames[13][3][10] = 8'had;
frames[13][3][11] = 8'h89;
frames[13][3][12] = 8'h88;
frames[13][3][13] = 8'h89;
frames[13][3][14] = 8'h68;
frames[13][3][15] = 8'h64;
frames[13][3][16] = 8'hb1;
frames[13][3][17] = 8'hd5;
frames[13][3][18] = 8'hd5;
frames[13][3][19] = 8'hd5;
frames[13][3][20] = 8'hb1;
frames[13][3][21] = 8'h8d;
frames[13][3][22] = 8'h48;
frames[13][3][23] = 8'h20;
frames[13][3][24] = 8'h20;
frames[13][3][25] = 8'h24;
frames[13][3][26] = 8'h24;
frames[13][3][27] = 8'h69;
frames[13][3][28] = 8'h91;
frames[13][3][29] = 8'h69;
frames[13][3][30] = 8'h44;
frames[13][3][31] = 8'h48;
frames[13][3][32] = 8'h48;
frames[13][3][33] = 8'h48;
frames[13][3][34] = 8'h48;
frames[13][3][35] = 8'h48;
frames[13][3][36] = 8'h8d;
frames[13][3][37] = 8'h49;
frames[13][3][38] = 8'h49;
frames[13][3][39] = 8'h6e;
frames[13][4][0] = 8'hfa;
frames[13][4][1] = 8'hfa;
frames[13][4][2] = 8'hfa;
frames[13][4][3] = 8'hff;
frames[13][4][4] = 8'hff;
frames[13][4][5] = 8'hff;
frames[13][4][6] = 8'hfa;
frames[13][4][7] = 8'hd2;
frames[13][4][8] = 8'had;
frames[13][4][9] = 8'had;
frames[13][4][10] = 8'had;
frames[13][4][11] = 8'had;
frames[13][4][12] = 8'h88;
frames[13][4][13] = 8'h89;
frames[13][4][14] = 8'h89;
frames[13][4][15] = 8'h64;
frames[13][4][16] = 8'h8d;
frames[13][4][17] = 8'hb1;
frames[13][4][18] = 8'h8d;
frames[13][4][19] = 8'h69;
frames[13][4][20] = 8'h44;
frames[13][4][21] = 8'h24;
frames[13][4][22] = 8'h20;
frames[13][4][23] = 8'h24;
frames[13][4][24] = 8'h48;
frames[13][4][25] = 8'h8d;
frames[13][4][26] = 8'hb1;
frames[13][4][27] = 8'hb1;
frames[13][4][28] = 8'hb1;
frames[13][4][29] = 8'hb1;
frames[13][4][30] = 8'hb5;
frames[13][4][31] = 8'hb5;
frames[13][4][32] = 8'hb1;
frames[13][4][33] = 8'hb1;
frames[13][4][34] = 8'hb1;
frames[13][4][35] = 8'h8d;
frames[13][4][36] = 8'hb2;
frames[13][4][37] = 8'h91;
frames[13][4][38] = 8'h91;
frames[13][4][39] = 8'h6d;
frames[13][5][0] = 8'hfa;
frames[13][5][1] = 8'hfa;
frames[13][5][2] = 8'hff;
frames[13][5][3] = 8'hff;
frames[13][5][4] = 8'hff;
frames[13][5][5] = 8'hff;
frames[13][5][6] = 8'hfb;
frames[13][5][7] = 8'hfa;
frames[13][5][8] = 8'had;
frames[13][5][9] = 8'had;
frames[13][5][10] = 8'h89;
frames[13][5][11] = 8'had;
frames[13][5][12] = 8'h89;
frames[13][5][13] = 8'h68;
frames[13][5][14] = 8'h89;
frames[13][5][15] = 8'h88;
frames[13][5][16] = 8'h68;
frames[13][5][17] = 8'h44;
frames[13][5][18] = 8'h24;
frames[13][5][19] = 8'h24;
frames[13][5][20] = 8'h24;
frames[13][5][21] = 8'h24;
frames[13][5][22] = 8'h24;
frames[13][5][23] = 8'h6d;
frames[13][5][24] = 8'hb1;
frames[13][5][25] = 8'hb1;
frames[13][5][26] = 8'hb1;
frames[13][5][27] = 8'hb1;
frames[13][5][28] = 8'hb1;
frames[13][5][29] = 8'hb1;
frames[13][5][30] = 8'hb5;
frames[13][5][31] = 8'hb5;
frames[13][5][32] = 8'hb5;
frames[13][5][33] = 8'hb1;
frames[13][5][34] = 8'hb1;
frames[13][5][35] = 8'hb1;
frames[13][5][36] = 8'h8d;
frames[13][5][37] = 8'hd6;
frames[13][5][38] = 8'hb2;
frames[13][5][39] = 8'h6d;
frames[13][6][0] = 8'hfa;
frames[13][6][1] = 8'hff;
frames[13][6][2] = 8'hff;
frames[13][6][3] = 8'hff;
frames[13][6][4] = 8'hff;
frames[13][6][5] = 8'hfe;
frames[13][6][6] = 8'hfb;
frames[13][6][7] = 8'hfa;
frames[13][6][8] = 8'hd6;
frames[13][6][9] = 8'had;
frames[13][6][10] = 8'h89;
frames[13][6][11] = 8'ha9;
frames[13][6][12] = 8'had;
frames[13][6][13] = 8'h64;
frames[13][6][14] = 8'h64;
frames[13][6][15] = 8'h88;
frames[13][6][16] = 8'h68;
frames[13][6][17] = 8'h44;
frames[13][6][18] = 8'h24;
frames[13][6][19] = 8'h24;
frames[13][6][20] = 8'h24;
frames[13][6][21] = 8'h49;
frames[13][6][22] = 8'hb1;
frames[13][6][23] = 8'hb2;
frames[13][6][24] = 8'hb1;
frames[13][6][25] = 8'h91;
frames[13][6][26] = 8'hb1;
frames[13][6][27] = 8'hb1;
frames[13][6][28] = 8'hd5;
frames[13][6][29] = 8'hd5;
frames[13][6][30] = 8'hd5;
frames[13][6][31] = 8'hd5;
frames[13][6][32] = 8'hb5;
frames[13][6][33] = 8'hb1;
frames[13][6][34] = 8'hb1;
frames[13][6][35] = 8'h8d;
frames[13][6][36] = 8'h8d;
frames[13][6][37] = 8'hb1;
frames[13][6][38] = 8'h8d;
frames[13][6][39] = 8'h68;
frames[13][7][0] = 8'hfa;
frames[13][7][1] = 8'hfe;
frames[13][7][2] = 8'hff;
frames[13][7][3] = 8'hfa;
frames[13][7][4] = 8'hfa;
frames[13][7][5] = 8'hfa;
frames[13][7][6] = 8'hfb;
frames[13][7][7] = 8'hff;
frames[13][7][8] = 8'hfa;
frames[13][7][9] = 8'hb1;
frames[13][7][10] = 8'had;
frames[13][7][11] = 8'h89;
frames[13][7][12] = 8'had;
frames[13][7][13] = 8'h88;
frames[13][7][14] = 8'h64;
frames[13][7][15] = 8'h88;
frames[13][7][16] = 8'h68;
frames[13][7][17] = 8'h44;
frames[13][7][18] = 8'h24;
frames[13][7][19] = 8'h48;
frames[13][7][20] = 8'hb1;
frames[13][7][21] = 8'hd6;
frames[13][7][22] = 8'hb1;
frames[13][7][23] = 8'hb1;
frames[13][7][24] = 8'hb1;
frames[13][7][25] = 8'hb1;
frames[13][7][26] = 8'hb1;
frames[13][7][27] = 8'hb5;
frames[13][7][28] = 8'hd5;
frames[13][7][29] = 8'hd6;
frames[13][7][30] = 8'hda;
frames[13][7][31] = 8'hd6;
frames[13][7][32] = 8'hd6;
frames[13][7][33] = 8'hb1;
frames[13][7][34] = 8'hb1;
frames[13][7][35] = 8'h8d;
frames[13][7][36] = 8'h91;
frames[13][7][37] = 8'hb1;
frames[13][7][38] = 8'hb1;
frames[13][7][39] = 8'h68;
frames[13][8][0] = 8'hfa;
frames[13][8][1] = 8'hff;
frames[13][8][2] = 8'hfb;
frames[13][8][3] = 8'hff;
frames[13][8][4] = 8'hff;
frames[13][8][5] = 8'hff;
frames[13][8][6] = 8'hfb;
frames[13][8][7] = 8'hb6;
frames[13][8][8] = 8'h8d;
frames[13][8][9] = 8'h69;
frames[13][8][10] = 8'had;
frames[13][8][11] = 8'had;
frames[13][8][12] = 8'had;
frames[13][8][13] = 8'had;
frames[13][8][14] = 8'h88;
frames[13][8][15] = 8'h64;
frames[13][8][16] = 8'h48;
frames[13][8][17] = 8'h69;
frames[13][8][18] = 8'h91;
frames[13][8][19] = 8'hb6;
frames[13][8][20] = 8'hd6;
frames[13][8][21] = 8'hb1;
frames[13][8][22] = 8'hb1;
frames[13][8][23] = 8'hb1;
frames[13][8][24] = 8'hb1;
frames[13][8][25] = 8'hd5;
frames[13][8][26] = 8'hb1;
frames[13][8][27] = 8'hd5;
frames[13][8][28] = 8'hd6;
frames[13][8][29] = 8'hd6;
frames[13][8][30] = 8'hd6;
frames[13][8][31] = 8'hb5;
frames[13][8][32] = 8'hb5;
frames[13][8][33] = 8'h91;
frames[13][8][34] = 8'hb1;
frames[13][8][35] = 8'hb5;
frames[13][8][36] = 8'hb1;
frames[13][8][37] = 8'hb1;
frames[13][8][38] = 8'hb1;
frames[13][8][39] = 8'h8d;
frames[13][9][0] = 8'hff;
frames[13][9][1] = 8'hff;
frames[13][9][2] = 8'hff;
frames[13][9][3] = 8'hff;
frames[13][9][4] = 8'hd6;
frames[13][9][5] = 8'h8d;
frames[13][9][6] = 8'h49;
frames[13][9][7] = 8'h24;
frames[13][9][8] = 8'h24;
frames[13][9][9] = 8'h44;
frames[13][9][10] = 8'ha9;
frames[13][9][11] = 8'h88;
frames[13][9][12] = 8'hb1;
frames[13][9][13] = 8'hd1;
frames[13][9][14] = 8'had;
frames[13][9][15] = 8'h89;
frames[13][9][16] = 8'hb2;
frames[13][9][17] = 8'hb6;
frames[13][9][18] = 8'hb6;
frames[13][9][19] = 8'hb6;
frames[13][9][20] = 8'hb1;
frames[13][9][21] = 8'hb1;
frames[13][9][22] = 8'hb1;
frames[13][9][23] = 8'hb1;
frames[13][9][24] = 8'hb1;
frames[13][9][25] = 8'hb1;
frames[13][9][26] = 8'hb1;
frames[13][9][27] = 8'hb1;
frames[13][9][28] = 8'hd5;
frames[13][9][29] = 8'hb5;
frames[13][9][30] = 8'hb5;
frames[13][9][31] = 8'hb1;
frames[13][9][32] = 8'h8d;
frames[13][9][33] = 8'h68;
frames[13][9][34] = 8'h68;
frames[13][9][35] = 8'hb1;
frames[13][9][36] = 8'hb1;
frames[13][9][37] = 8'hb1;
frames[13][9][38] = 8'hb1;
frames[13][9][39] = 8'h8d;
frames[13][10][0] = 8'hfb;
frames[13][10][1] = 8'hda;
frames[13][10][2] = 8'h92;
frames[13][10][3] = 8'h49;
frames[13][10][4] = 8'h24;
frames[13][10][5] = 8'h24;
frames[13][10][6] = 8'h24;
frames[13][10][7] = 8'h24;
frames[13][10][8] = 8'h24;
frames[13][10][9] = 8'h24;
frames[13][10][10] = 8'h88;
frames[13][10][11] = 8'h89;
frames[13][10][12] = 8'had;
frames[13][10][13] = 8'hd5;
frames[13][10][14] = 8'hb1;
frames[13][10][15] = 8'hb1;
frames[13][10][16] = 8'hb6;
frames[13][10][17] = 8'hb6;
frames[13][10][18] = 8'hb5;
frames[13][10][19] = 8'hb1;
frames[13][10][20] = 8'hb1;
frames[13][10][21] = 8'h8d;
frames[13][10][22] = 8'h8d;
frames[13][10][23] = 8'hb1;
frames[13][10][24] = 8'hb1;
frames[13][10][25] = 8'h8d;
frames[13][10][26] = 8'h8d;
frames[13][10][27] = 8'h8d;
frames[13][10][28] = 8'hb1;
frames[13][10][29] = 8'h91;
frames[13][10][30] = 8'hb1;
frames[13][10][31] = 8'hb1;
frames[13][10][32] = 8'h91;
frames[13][10][33] = 8'h91;
frames[13][10][34] = 8'h91;
frames[13][10][35] = 8'hd6;
frames[13][10][36] = 8'hb2;
frames[13][10][37] = 8'h8d;
frames[13][10][38] = 8'h48;
frames[13][10][39] = 8'h48;
frames[13][11][0] = 8'h69;
frames[13][11][1] = 8'h44;
frames[13][11][2] = 8'h24;
frames[13][11][3] = 8'h24;
frames[13][11][4] = 8'h24;
frames[13][11][5] = 8'h48;
frames[13][11][6] = 8'h44;
frames[13][11][7] = 8'h44;
frames[13][11][8] = 8'h68;
frames[13][11][9] = 8'h6d;
frames[13][11][10] = 8'hb1;
frames[13][11][11] = 8'h8d;
frames[13][11][12] = 8'h8d;
frames[13][11][13] = 8'hd1;
frames[13][11][14] = 8'hb1;
frames[13][11][15] = 8'hb6;
frames[13][11][16] = 8'hd6;
frames[13][11][17] = 8'hd6;
frames[13][11][18] = 8'h91;
frames[13][11][19] = 8'h8d;
frames[13][11][20] = 8'hb1;
frames[13][11][21] = 8'h91;
frames[13][11][22] = 8'hb1;
frames[13][11][23] = 8'hb1;
frames[13][11][24] = 8'hb1;
frames[13][11][25] = 8'h8d;
frames[13][11][26] = 8'h8d;
frames[13][11][27] = 8'h8d;
frames[13][11][28] = 8'hb1;
frames[13][11][29] = 8'hb5;
frames[13][11][30] = 8'hb1;
frames[13][11][31] = 8'hb1;
frames[13][11][32] = 8'hb1;
frames[13][11][33] = 8'h8d;
frames[13][11][34] = 8'h6d;
frames[13][11][35] = 8'h91;
frames[13][11][36] = 8'h8d;
frames[13][11][37] = 8'h44;
frames[13][11][38] = 8'h44;
frames[13][11][39] = 8'h44;
frames[13][12][0] = 8'h24;
frames[13][12][1] = 8'h24;
frames[13][12][2] = 8'h44;
frames[13][12][3] = 8'h44;
frames[13][12][4] = 8'h8d;
frames[13][12][5] = 8'hb1;
frames[13][12][6] = 8'h88;
frames[13][12][7] = 8'h89;
frames[13][12][8] = 8'hd1;
frames[13][12][9] = 8'hd5;
frames[13][12][10] = 8'hd5;
frames[13][12][11] = 8'hb1;
frames[13][12][12] = 8'hb1;
frames[13][12][13] = 8'hd1;
frames[13][12][14] = 8'hb1;
frames[13][12][15] = 8'h68;
frames[13][12][16] = 8'h8d;
frames[13][12][17] = 8'hd2;
frames[13][12][18] = 8'h8d;
frames[13][12][19] = 8'h24;
frames[13][12][20] = 8'h24;
frames[13][12][21] = 8'h48;
frames[13][12][22] = 8'h8d;
frames[13][12][23] = 8'h8d;
frames[13][12][24] = 8'h6d;
frames[13][12][25] = 8'h8d;
frames[13][12][26] = 8'h68;
frames[13][12][27] = 8'h6d;
frames[13][12][28] = 8'h8d;
frames[13][12][29] = 8'h6d;
frames[13][12][30] = 8'h69;
frames[13][12][31] = 8'h68;
frames[13][12][32] = 8'h44;
frames[13][12][33] = 8'h44;
frames[13][12][34] = 8'h44;
frames[13][12][35] = 8'h8d;
frames[13][12][36] = 8'hb2;
frames[13][12][37] = 8'h48;
frames[13][12][38] = 8'h44;
frames[13][12][39] = 8'h44;
frames[13][13][0] = 8'h69;
frames[13][13][1] = 8'h69;
frames[13][13][2] = 8'had;
frames[13][13][3] = 8'hd1;
frames[13][13][4] = 8'hd1;
frames[13][13][5] = 8'hd1;
frames[13][13][6] = 8'had;
frames[13][13][7] = 8'hb1;
frames[13][13][8] = 8'hd5;
frames[13][13][9] = 8'hd6;
frames[13][13][10] = 8'hd5;
frames[13][13][11] = 8'hb1;
frames[13][13][12] = 8'hd1;
frames[13][13][13] = 8'hd5;
frames[13][13][14] = 8'hb1;
frames[13][13][15] = 8'h8c;
frames[13][13][16] = 8'h64;
frames[13][13][17] = 8'h8d;
frames[13][13][18] = 8'hb2;
frames[13][13][19] = 8'h6d;
frames[13][13][20] = 8'h24;
frames[13][13][21] = 8'h44;
frames[13][13][22] = 8'h8d;
frames[13][13][23] = 8'h6d;
frames[13][13][24] = 8'h69;
frames[13][13][25] = 8'h6d;
frames[13][13][26] = 8'h6d;
frames[13][13][27] = 8'h6d;
frames[13][13][28] = 8'h6d;
frames[13][13][29] = 8'h6d;
frames[13][13][30] = 8'h6d;
frames[13][13][31] = 8'h6d;
frames[13][13][32] = 8'h6d;
frames[13][13][33] = 8'h6d;
frames[13][13][34] = 8'h6d;
frames[13][13][35] = 8'h91;
frames[13][13][36] = 8'hb6;
frames[13][13][37] = 8'h6d;
frames[13][13][38] = 8'h68;
frames[13][13][39] = 8'h48;
frames[13][14][0] = 8'hd6;
frames[13][14][1] = 8'hd6;
frames[13][14][2] = 8'hb1;
frames[13][14][3] = 8'had;
frames[13][14][4] = 8'hd6;
frames[13][14][5] = 8'hd6;
frames[13][14][6] = 8'hb1;
frames[13][14][7] = 8'hb1;
frames[13][14][8] = 8'hd5;
frames[13][14][9] = 8'hd6;
frames[13][14][10] = 8'hd5;
frames[13][14][11] = 8'hb1;
frames[13][14][12] = 8'hb1;
frames[13][14][13] = 8'hb1;
frames[13][14][14] = 8'hb1;
frames[13][14][15] = 8'hb1;
frames[13][14][16] = 8'h68;
frames[13][14][17] = 8'h89;
frames[13][14][18] = 8'hb6;
frames[13][14][19] = 8'hd6;
frames[13][14][20] = 8'hb1;
frames[13][14][21] = 8'h91;
frames[13][14][22] = 8'hb6;
frames[13][14][23] = 8'hb6;
frames[13][14][24] = 8'hb2;
frames[13][14][25] = 8'hb2;
frames[13][14][26] = 8'hb2;
frames[13][14][27] = 8'h91;
frames[13][14][28] = 8'h8d;
frames[13][14][29] = 8'h8d;
frames[13][14][30] = 8'h8d;
frames[13][14][31] = 8'h8d;
frames[13][14][32] = 8'h8d;
frames[13][14][33] = 8'h6d;
frames[13][14][34] = 8'h6d;
frames[13][14][35] = 8'h8d;
frames[13][14][36] = 8'hb6;
frames[13][14][37] = 8'h6d;
frames[13][14][38] = 8'h6d;
frames[13][14][39] = 8'h6d;
frames[13][15][0] = 8'hda;
frames[13][15][1] = 8'hd6;
frames[13][15][2] = 8'hb1;
frames[13][15][3] = 8'hd6;
frames[13][15][4] = 8'hb1;
frames[13][15][5] = 8'hb1;
frames[13][15][6] = 8'hb1;
frames[13][15][7] = 8'hb1;
frames[13][15][8] = 8'hd6;
frames[13][15][9] = 8'hd6;
frames[13][15][10] = 8'hd5;
frames[13][15][11] = 8'hb1;
frames[13][15][12] = 8'hb1;
frames[13][15][13] = 8'hb1;
frames[13][15][14] = 8'had;
frames[13][15][15] = 8'h8d;
frames[13][15][16] = 8'h8d;
frames[13][15][17] = 8'had;
frames[13][15][18] = 8'hb1;
frames[13][15][19] = 8'hb1;
frames[13][15][20] = 8'h8d;
frames[13][15][21] = 8'hb1;
frames[13][15][22] = 8'hb6;
frames[13][15][23] = 8'hb2;
frames[13][15][24] = 8'hb2;
frames[13][15][25] = 8'h91;
frames[13][15][26] = 8'h8d;
frames[13][15][27] = 8'h8d;
frames[13][15][28] = 8'h8d;
frames[13][15][29] = 8'h8d;
frames[13][15][30] = 8'h8d;
frames[13][15][31] = 8'h8d;
frames[13][15][32] = 8'h69;
frames[13][15][33] = 8'h44;
frames[13][15][34] = 8'h24;
frames[13][15][35] = 8'hb6;
frames[13][15][36] = 8'hff;
frames[13][15][37] = 8'h69;
frames[13][15][38] = 8'h44;
frames[13][15][39] = 8'h44;
frames[13][16][0] = 8'hd5;
frames[13][16][1] = 8'hd5;
frames[13][16][2] = 8'hd6;
frames[13][16][3] = 8'hb5;
frames[13][16][4] = 8'had;
frames[13][16][5] = 8'h8d;
frames[13][16][6] = 8'hd5;
frames[13][16][7] = 8'hb1;
frames[13][16][8] = 8'hb1;
frames[13][16][9] = 8'hb1;
frames[13][16][10] = 8'hb1;
frames[13][16][11] = 8'h8d;
frames[13][16][12] = 8'hb1;
frames[13][16][13] = 8'hb1;
frames[13][16][14] = 8'had;
frames[13][16][15] = 8'h64;
frames[13][16][16] = 8'h89;
frames[13][16][17] = 8'h89;
frames[13][16][18] = 8'hb1;
frames[13][16][19] = 8'hb1;
frames[13][16][20] = 8'hb1;
frames[13][16][21] = 8'hb1;
frames[13][16][22] = 8'hb2;
frames[13][16][23] = 8'h91;
frames[13][16][24] = 8'h91;
frames[13][16][25] = 8'hb2;
frames[13][16][26] = 8'hb6;
frames[13][16][27] = 8'hb2;
frames[13][16][28] = 8'h92;
frames[13][16][29] = 8'h8d;
frames[13][16][30] = 8'h69;
frames[13][16][31] = 8'h48;
frames[13][16][32] = 8'h24;
frames[13][16][33] = 8'h24;
frames[13][16][34] = 8'h24;
frames[13][16][35] = 8'h6d;
frames[13][16][36] = 8'hb6;
frames[13][16][37] = 8'h49;
frames[13][16][38] = 8'h44;
frames[13][16][39] = 8'h44;
frames[13][17][0] = 8'hd5;
frames[13][17][1] = 8'hb1;
frames[13][17][2] = 8'hb1;
frames[13][17][3] = 8'had;
frames[13][17][4] = 8'h8d;
frames[13][17][5] = 8'h8c;
frames[13][17][6] = 8'hb1;
frames[13][17][7] = 8'hd6;
frames[13][17][8] = 8'h88;
frames[13][17][9] = 8'had;
frames[13][17][10] = 8'hb1;
frames[13][17][11] = 8'h8d;
frames[13][17][12] = 8'hb1;
frames[13][17][13] = 8'hb1;
frames[13][17][14] = 8'had;
frames[13][17][15] = 8'h8d;
frames[13][17][16] = 8'h88;
frames[13][17][17] = 8'h89;
frames[13][17][18] = 8'hb1;
frames[13][17][19] = 8'hb1;
frames[13][17][20] = 8'h8d;
frames[13][17][21] = 8'hb2;
frames[13][17][22] = 8'hb2;
frames[13][17][23] = 8'hb6;
frames[13][17][24] = 8'hb6;
frames[13][17][25] = 8'hb6;
frames[13][17][26] = 8'hd6;
frames[13][17][27] = 8'hb2;
frames[13][17][28] = 8'h69;
frames[13][17][29] = 8'h44;
frames[13][17][30] = 8'h24;
frames[13][17][31] = 8'h24;
frames[13][17][32] = 8'h24;
frames[13][17][33] = 8'h24;
frames[13][17][34] = 8'h44;
frames[13][17][35] = 8'h44;
frames[13][17][36] = 8'h44;
frames[13][17][37] = 8'h44;
frames[13][17][38] = 8'h44;
frames[13][17][39] = 8'h44;
frames[13][18][0] = 8'had;
frames[13][18][1] = 8'h88;
frames[13][18][2] = 8'h8c;
frames[13][18][3] = 8'hd1;
frames[13][18][4] = 8'hd6;
frames[13][18][5] = 8'hb1;
frames[13][18][6] = 8'hb1;
frames[13][18][7] = 8'hb1;
frames[13][18][8] = 8'had;
frames[13][18][9] = 8'h88;
frames[13][18][10] = 8'h88;
frames[13][18][11] = 8'had;
frames[13][18][12] = 8'hd5;
frames[13][18][13] = 8'hb1;
frames[13][18][14] = 8'h8d;
frames[13][18][15] = 8'hb1;
frames[13][18][16] = 8'h89;
frames[13][18][17] = 8'h89;
frames[13][18][18] = 8'h91;
frames[13][18][19] = 8'h69;
frames[13][18][20] = 8'h6d;
frames[13][18][21] = 8'h8d;
frames[13][18][22] = 8'hb6;
frames[13][18][23] = 8'hd6;
frames[13][18][24] = 8'hb6;
frames[13][18][25] = 8'h91;
frames[13][18][26] = 8'h8d;
frames[13][18][27] = 8'h69;
frames[13][18][28] = 8'h24;
frames[13][18][29] = 8'h24;
frames[13][18][30] = 8'h24;
frames[13][18][31] = 8'h24;
frames[13][18][32] = 8'h44;
frames[13][18][33] = 8'h44;
frames[13][18][34] = 8'h48;
frames[13][18][35] = 8'h69;
frames[13][18][36] = 8'h6d;
frames[13][18][37] = 8'h68;
frames[13][18][38] = 8'h68;
frames[13][18][39] = 8'h8d;
frames[13][19][0] = 8'hb1;
frames[13][19][1] = 8'hb1;
frames[13][19][2] = 8'hd6;
frames[13][19][3] = 8'hb5;
frames[13][19][4] = 8'hd5;
frames[13][19][5] = 8'hd6;
frames[13][19][6] = 8'hd6;
frames[13][19][7] = 8'hb1;
frames[13][19][8] = 8'hb1;
frames[13][19][9] = 8'h88;
frames[13][19][10] = 8'h88;
frames[13][19][11] = 8'h89;
frames[13][19][12] = 8'hb1;
frames[13][19][13] = 8'hb1;
frames[13][19][14] = 8'hb1;
frames[13][19][15] = 8'hb1;
frames[13][19][16] = 8'h8d;
frames[13][19][17] = 8'h68;
frames[13][19][18] = 8'h69;
frames[13][19][19] = 8'hb2;
frames[13][19][20] = 8'hb1;
frames[13][19][21] = 8'h68;
frames[13][19][22] = 8'h8d;
frames[13][19][23] = 8'h91;
frames[13][19][24] = 8'h91;
frames[13][19][25] = 8'h8d;
frames[13][19][26] = 8'h6d;
frames[13][19][27] = 8'h69;
frames[13][19][28] = 8'h6d;
frames[13][19][29] = 8'h69;
frames[13][19][30] = 8'h68;
frames[13][19][31] = 8'h68;
frames[13][19][32] = 8'h68;
frames[13][19][33] = 8'h68;
frames[13][19][34] = 8'h6d;
frames[13][19][35] = 8'h8d;
frames[13][19][36] = 8'h8d;
frames[13][19][37] = 8'h8d;
frames[13][19][38] = 8'h8d;
frames[13][19][39] = 8'h8d;
frames[13][20][0] = 8'h91;
frames[13][20][1] = 8'hb1;
frames[13][20][2] = 8'hb5;
frames[13][20][3] = 8'hb1;
frames[13][20][4] = 8'hb1;
frames[13][20][5] = 8'hb5;
frames[13][20][6] = 8'hd6;
frames[13][20][7] = 8'hd6;
frames[13][20][8] = 8'hd6;
frames[13][20][9] = 8'hb1;
frames[13][20][10] = 8'hb5;
frames[13][20][11] = 8'hb1;
frames[13][20][12] = 8'hb1;
frames[13][20][13] = 8'hb1;
frames[13][20][14] = 8'hb2;
frames[13][20][15] = 8'h68;
frames[13][20][16] = 8'h24;
frames[13][20][17] = 8'h69;
frames[13][20][18] = 8'hb6;
frames[13][20][19] = 8'hb6;
frames[13][20][20] = 8'h8d;
frames[13][20][21] = 8'h69;
frames[13][20][22] = 8'h68;
frames[13][20][23] = 8'h68;
frames[13][20][24] = 8'h68;
frames[13][20][25] = 8'h69;
frames[13][20][26] = 8'h68;
frames[13][20][27] = 8'h8d;
frames[13][20][28] = 8'h91;
frames[13][20][29] = 8'hd6;
frames[13][20][30] = 8'hb1;
frames[13][20][31] = 8'h8d;
frames[13][20][32] = 8'h8d;
frames[13][20][33] = 8'h8d;
frames[13][20][34] = 8'hb1;
frames[13][20][35] = 8'hb1;
frames[13][20][36] = 8'hb1;
frames[13][20][37] = 8'hb1;
frames[13][20][38] = 8'hb1;
frames[13][20][39] = 8'hb1;
frames[13][21][0] = 8'h44;
frames[13][21][1] = 8'h68;
frames[13][21][2] = 8'h8d;
frames[13][21][3] = 8'h91;
frames[13][21][4] = 8'hb1;
frames[13][21][5] = 8'hb1;
frames[13][21][6] = 8'hb1;
frames[13][21][7] = 8'hb1;
frames[13][21][8] = 8'hb1;
frames[13][21][9] = 8'hb1;
frames[13][21][10] = 8'h8d;
frames[13][21][11] = 8'h8d;
frames[13][21][12] = 8'h69;
frames[13][21][13] = 8'h68;
frames[13][21][14] = 8'h6d;
frames[13][21][15] = 8'h24;
frames[13][21][16] = 8'h44;
frames[13][21][17] = 8'h69;
frames[13][21][18] = 8'h49;
frames[13][21][19] = 8'h24;
frames[13][21][20] = 8'h24;
frames[13][21][21] = 8'h68;
frames[13][21][22] = 8'h69;
frames[13][21][23] = 8'h69;
frames[13][21][24] = 8'h8d;
frames[13][21][25] = 8'hb1;
frames[13][21][26] = 8'h91;
frames[13][21][27] = 8'hb1;
frames[13][21][28] = 8'hb1;
frames[13][21][29] = 8'hd6;
frames[13][21][30] = 8'hd6;
frames[13][21][31] = 8'hd6;
frames[13][21][32] = 8'hd6;
frames[13][21][33] = 8'hd5;
frames[13][21][34] = 8'hd6;
frames[13][21][35] = 8'hd6;
frames[13][21][36] = 8'hd1;
frames[13][21][37] = 8'hd5;
frames[13][21][38] = 8'hd5;
frames[13][21][39] = 8'hb1;
frames[13][22][0] = 8'hb2;
frames[13][22][1] = 8'h69;
frames[13][22][2] = 8'h20;
frames[13][22][3] = 8'h20;
frames[13][22][4] = 8'h24;
frames[13][22][5] = 8'h24;
frames[13][22][6] = 8'h24;
frames[13][22][7] = 8'h24;
frames[13][22][8] = 8'h24;
frames[13][22][9] = 8'h24;
frames[13][22][10] = 8'h24;
frames[13][22][11] = 8'h24;
frames[13][22][12] = 8'h24;
frames[13][22][13] = 8'h44;
frames[13][22][14] = 8'h24;
frames[13][22][15] = 8'h24;
frames[13][22][16] = 8'h24;
frames[13][22][17] = 8'h24;
frames[13][22][18] = 8'h20;
frames[13][22][19] = 8'h20;
frames[13][22][20] = 8'h20;
frames[13][22][21] = 8'h44;
frames[13][22][22] = 8'h69;
frames[13][22][23] = 8'h8d;
frames[13][22][24] = 8'hb1;
frames[13][22][25] = 8'hd6;
frames[13][22][26] = 8'hd6;
frames[13][22][27] = 8'hb6;
frames[13][22][28] = 8'hb6;
frames[13][22][29] = 8'hd6;
frames[13][22][30] = 8'hd6;
frames[13][22][31] = 8'hd6;
frames[13][22][32] = 8'hd5;
frames[13][22][33] = 8'hd5;
frames[13][22][34] = 8'hd5;
frames[13][22][35] = 8'hd5;
frames[13][22][36] = 8'hb5;
frames[13][22][37] = 8'hb1;
frames[13][22][38] = 8'hb1;
frames[13][22][39] = 8'hb1;
frames[13][23][0] = 8'hd6;
frames[13][23][1] = 8'hfb;
frames[13][23][2] = 8'hd6;
frames[13][23][3] = 8'h6d;
frames[13][23][4] = 8'h24;
frames[13][23][5] = 8'h24;
frames[13][23][6] = 8'h44;
frames[13][23][7] = 8'h69;
frames[13][23][8] = 8'h6d;
frames[13][23][9] = 8'h6d;
frames[13][23][10] = 8'h69;
frames[13][23][11] = 8'h49;
frames[13][23][12] = 8'h44;
frames[13][23][13] = 8'h44;
frames[13][23][14] = 8'h24;
frames[13][23][15] = 8'h24;
frames[13][23][16] = 8'h24;
frames[13][23][17] = 8'h20;
frames[13][23][18] = 8'h20;
frames[13][23][19] = 8'h24;
frames[13][23][20] = 8'h20;
frames[13][23][21] = 8'h44;
frames[13][23][22] = 8'h68;
frames[13][23][23] = 8'h8d;
frames[13][23][24] = 8'h8d;
frames[13][23][25] = 8'h8d;
frames[13][23][26] = 8'hb1;
frames[13][23][27] = 8'hb1;
frames[13][23][28] = 8'hb1;
frames[13][23][29] = 8'hb1;
frames[13][23][30] = 8'hb1;
frames[13][23][31] = 8'hb1;
frames[13][23][32] = 8'hb1;
frames[13][23][33] = 8'hb1;
frames[13][23][34] = 8'hb1;
frames[13][23][35] = 8'hb1;
frames[13][23][36] = 8'hb1;
frames[13][23][37] = 8'hb1;
frames[13][23][38] = 8'hb1;
frames[13][23][39] = 8'hb5;
frames[13][24][0] = 8'h44;
frames[13][24][1] = 8'h69;
frames[13][24][2] = 8'h92;
frames[13][24][3] = 8'hd6;
frames[13][24][4] = 8'hda;
frames[13][24][5] = 8'hdb;
frames[13][24][6] = 8'hfb;
frames[13][24][7] = 8'hfb;
frames[13][24][8] = 8'hdb;
frames[13][24][9] = 8'hb2;
frames[13][24][10] = 8'h69;
frames[13][24][11] = 8'h44;
frames[13][24][12] = 8'h24;
frames[13][24][13] = 8'h24;
frames[13][24][14] = 8'h20;
frames[13][24][15] = 8'h20;
frames[13][24][16] = 8'h20;
frames[13][24][17] = 8'h20;
frames[13][24][18] = 8'h24;
frames[13][24][19] = 8'h44;
frames[13][24][20] = 8'h44;
frames[13][24][21] = 8'h44;
frames[13][24][22] = 8'h68;
frames[13][24][23] = 8'h8d;
frames[13][24][24] = 8'hd6;
frames[13][24][25] = 8'hd6;
frames[13][24][26] = 8'hb5;
frames[13][24][27] = 8'hb5;
frames[13][24][28] = 8'hb5;
frames[13][24][29] = 8'hb5;
frames[13][24][30] = 8'hb5;
frames[13][24][31] = 8'hb1;
frames[13][24][32] = 8'hb5;
frames[13][24][33] = 8'hb1;
frames[13][24][34] = 8'hb1;
frames[13][24][35] = 8'hd5;
frames[13][24][36] = 8'hb5;
frames[13][24][37] = 8'hd5;
frames[13][24][38] = 8'hd6;
frames[13][24][39] = 8'hd6;
frames[13][25][0] = 8'h44;
frames[13][25][1] = 8'h44;
frames[13][25][2] = 8'h24;
frames[13][25][3] = 8'h44;
frames[13][25][4] = 8'h49;
frames[13][25][5] = 8'h8d;
frames[13][25][6] = 8'hb6;
frames[13][25][7] = 8'hb6;
frames[13][25][8] = 8'h92;
frames[13][25][9] = 8'h48;
frames[13][25][10] = 8'h24;
frames[13][25][11] = 8'h24;
frames[13][25][12] = 8'h20;
frames[13][25][13] = 8'h20;
frames[13][25][14] = 8'h24;
frames[13][25][15] = 8'h24;
frames[13][25][16] = 8'h24;
frames[13][25][17] = 8'h44;
frames[13][25][18] = 8'h44;
frames[13][25][19] = 8'h44;
frames[13][25][20] = 8'h64;
frames[13][25][21] = 8'h68;
frames[13][25][22] = 8'h88;
frames[13][25][23] = 8'h8d;
frames[13][25][24] = 8'hfa;
frames[13][25][25] = 8'hff;
frames[13][25][26] = 8'hd6;
frames[13][25][27] = 8'hb5;
frames[13][25][28] = 8'hb5;
frames[13][25][29] = 8'hd5;
frames[13][25][30] = 8'hd5;
frames[13][25][31] = 8'hb5;
frames[13][25][32] = 8'hb5;
frames[13][25][33] = 8'hd5;
frames[13][25][34] = 8'hb5;
frames[13][25][35] = 8'hd5;
frames[13][25][36] = 8'hd5;
frames[13][25][37] = 8'hd5;
frames[13][25][38] = 8'hd6;
frames[13][25][39] = 8'hd6;
frames[13][26][0] = 8'h44;
frames[13][26][1] = 8'h24;
frames[13][26][2] = 8'h24;
frames[13][26][3] = 8'h24;
frames[13][26][4] = 8'h24;
frames[13][26][5] = 8'h24;
frames[13][26][6] = 8'h24;
frames[13][26][7] = 8'h44;
frames[13][26][8] = 8'h24;
frames[13][26][9] = 8'h00;
frames[13][26][10] = 8'h20;
frames[13][26][11] = 8'h24;
frames[13][26][12] = 8'h20;
frames[13][26][13] = 8'h20;
frames[13][26][14] = 8'h44;
frames[13][26][15] = 8'h44;
frames[13][26][16] = 8'h44;
frames[13][26][17] = 8'h44;
frames[13][26][18] = 8'h68;
frames[13][26][19] = 8'h68;
frames[13][26][20] = 8'h68;
frames[13][26][21] = 8'h8c;
frames[13][26][22] = 8'had;
frames[13][26][23] = 8'had;
frames[13][26][24] = 8'hb1;
frames[13][26][25] = 8'hd6;
frames[13][26][26] = 8'hd6;
frames[13][26][27] = 8'hb5;
frames[13][26][28] = 8'hb5;
frames[13][26][29] = 8'hb1;
frames[13][26][30] = 8'hb5;
frames[13][26][31] = 8'hb5;
frames[13][26][32] = 8'hb5;
frames[13][26][33] = 8'hb5;
frames[13][26][34] = 8'hb5;
frames[13][26][35] = 8'hd6;
frames[13][26][36] = 8'hd6;
frames[13][26][37] = 8'hb6;
frames[13][26][38] = 8'hb5;
frames[13][26][39] = 8'hb5;
frames[13][27][0] = 8'h44;
frames[13][27][1] = 8'h44;
frames[13][27][2] = 8'h24;
frames[13][27][3] = 8'h24;
frames[13][27][4] = 8'h24;
frames[13][27][5] = 8'h24;
frames[13][27][6] = 8'h24;
frames[13][27][7] = 8'h44;
frames[13][27][8] = 8'h24;
frames[13][27][9] = 8'h20;
frames[13][27][10] = 8'h20;
frames[13][27][11] = 8'h24;
frames[13][27][12] = 8'h44;
frames[13][27][13] = 8'h44;
frames[13][27][14] = 8'h64;
frames[13][27][15] = 8'h68;
frames[13][27][16] = 8'h68;
frames[13][27][17] = 8'h68;
frames[13][27][18] = 8'h68;
frames[13][27][19] = 8'h68;
frames[13][27][20] = 8'h8c;
frames[13][27][21] = 8'had;
frames[13][27][22] = 8'hb1;
frames[13][27][23] = 8'hb1;
frames[13][27][24] = 8'hb1;
frames[13][27][25] = 8'hb1;
frames[13][27][26] = 8'hb5;
frames[13][27][27] = 8'hb5;
frames[13][27][28] = 8'hb5;
frames[13][27][29] = 8'hb1;
frames[13][27][30] = 8'hb1;
frames[13][27][31] = 8'hb5;
frames[13][27][32] = 8'hb5;
frames[13][27][33] = 8'hb1;
frames[13][27][34] = 8'hb1;
frames[13][27][35] = 8'hb5;
frames[13][27][36] = 8'hb5;
frames[13][27][37] = 8'hb1;
frames[13][27][38] = 8'hb1;
frames[13][27][39] = 8'hb1;
frames[13][28][0] = 8'h44;
frames[13][28][1] = 8'h44;
frames[13][28][2] = 8'h44;
frames[13][28][3] = 8'h44;
frames[13][28][4] = 8'h44;
frames[13][28][5] = 8'h44;
frames[13][28][6] = 8'h44;
frames[13][28][7] = 8'h44;
frames[13][28][8] = 8'h44;
frames[13][28][9] = 8'h44;
frames[13][28][10] = 8'h44;
frames[13][28][11] = 8'h44;
frames[13][28][12] = 8'h44;
frames[13][28][13] = 8'h68;
frames[13][28][14] = 8'h68;
frames[13][28][15] = 8'h68;
frames[13][28][16] = 8'h68;
frames[13][28][17] = 8'h68;
frames[13][28][18] = 8'h68;
frames[13][28][19] = 8'h88;
frames[13][28][20] = 8'h8d;
frames[13][28][21] = 8'had;
frames[13][28][22] = 8'hb1;
frames[13][28][23] = 8'hb1;
frames[13][28][24] = 8'hb1;
frames[13][28][25] = 8'hb1;
frames[13][28][26] = 8'hb1;
frames[13][28][27] = 8'hd5;
frames[13][28][28] = 8'hd6;
frames[13][28][29] = 8'hb1;
frames[13][28][30] = 8'hb1;
frames[13][28][31] = 8'hb5;
frames[13][28][32] = 8'hd5;
frames[13][28][33] = 8'hb5;
frames[13][28][34] = 8'hb6;
frames[13][28][35] = 8'hb1;
frames[13][28][36] = 8'hb1;
frames[13][28][37] = 8'hb1;
frames[13][28][38] = 8'h91;
frames[13][28][39] = 8'h91;
frames[13][29][0] = 8'h68;
frames[13][29][1] = 8'h64;
frames[13][29][2] = 8'h44;
frames[13][29][3] = 8'h44;
frames[13][29][4] = 8'h44;
frames[13][29][5] = 8'h44;
frames[13][29][6] = 8'h44;
frames[13][29][7] = 8'h44;
frames[13][29][8] = 8'h44;
frames[13][29][9] = 8'h44;
frames[13][29][10] = 8'h44;
frames[13][29][11] = 8'h44;
frames[13][29][12] = 8'h68;
frames[13][29][13] = 8'h68;
frames[13][29][14] = 8'h68;
frames[13][29][15] = 8'h68;
frames[13][29][16] = 8'h68;
frames[13][29][17] = 8'h68;
frames[13][29][18] = 8'h88;
frames[13][29][19] = 8'h88;
frames[13][29][20] = 8'h8d;
frames[13][29][21] = 8'h8d;
frames[13][29][22] = 8'had;
frames[13][29][23] = 8'had;
frames[13][29][24] = 8'had;
frames[13][29][25] = 8'hb1;
frames[13][29][26] = 8'had;
frames[13][29][27] = 8'hb1;
frames[13][29][28] = 8'hd5;
frames[13][29][29] = 8'hb1;
frames[13][29][30] = 8'hb1;
frames[13][29][31] = 8'hb1;
frames[13][29][32] = 8'hb1;
frames[13][29][33] = 8'hb1;
frames[13][29][34] = 8'hb1;
frames[13][29][35] = 8'hb1;
frames[13][29][36] = 8'h91;
frames[13][29][37] = 8'h91;
frames[13][29][38] = 8'h8d;
frames[13][29][39] = 8'h8d;
frames[14][0][0] = 8'hd1;
frames[14][0][1] = 8'had;
frames[14][0][2] = 8'h8d;
frames[14][0][3] = 8'had;
frames[14][0][4] = 8'h89;
frames[14][0][5] = 8'h8d;
frames[14][0][6] = 8'h89;
frames[14][0][7] = 8'h44;
frames[14][0][8] = 8'h44;
frames[14][0][9] = 8'hb1;
frames[14][0][10] = 8'hd6;
frames[14][0][11] = 8'hd6;
frames[14][0][12] = 8'hd6;
frames[14][0][13] = 8'hd6;
frames[14][0][14] = 8'hd5;
frames[14][0][15] = 8'hd5;
frames[14][0][16] = 8'hd5;
frames[14][0][17] = 8'hd5;
frames[14][0][18] = 8'hd5;
frames[14][0][19] = 8'hd5;
frames[14][0][20] = 8'hd5;
frames[14][0][21] = 8'hd5;
frames[14][0][22] = 8'hd5;
frames[14][0][23] = 8'hd5;
frames[14][0][24] = 8'hd5;
frames[14][0][25] = 8'hd5;
frames[14][0][26] = 8'hd5;
frames[14][0][27] = 8'hb1;
frames[14][0][28] = 8'hb1;
frames[14][0][29] = 8'h69;
frames[14][0][30] = 8'h48;
frames[14][0][31] = 8'h44;
frames[14][0][32] = 8'h49;
frames[14][0][33] = 8'h6d;
frames[14][0][34] = 8'h8d;
frames[14][0][35] = 8'h91;
frames[14][0][36] = 8'h6d;
frames[14][0][37] = 8'h8d;
frames[14][0][38] = 8'h6d;
frames[14][0][39] = 8'h44;
frames[14][1][0] = 8'hd1;
frames[14][1][1] = 8'had;
frames[14][1][2] = 8'h89;
frames[14][1][3] = 8'had;
frames[14][1][4] = 8'h89;
frames[14][1][5] = 8'had;
frames[14][1][6] = 8'h89;
frames[14][1][7] = 8'h40;
frames[14][1][8] = 8'h68;
frames[14][1][9] = 8'hd6;
frames[14][1][10] = 8'hd6;
frames[14][1][11] = 8'hd6;
frames[14][1][12] = 8'hd6;
frames[14][1][13] = 8'hd6;
frames[14][1][14] = 8'hd5;
frames[14][1][15] = 8'hd5;
frames[14][1][16] = 8'hd5;
frames[14][1][17] = 8'hd5;
frames[14][1][18] = 8'hd5;
frames[14][1][19] = 8'hd5;
frames[14][1][20] = 8'hd6;
frames[14][1][21] = 8'hd6;
frames[14][1][22] = 8'hd5;
frames[14][1][23] = 8'hd5;
frames[14][1][24] = 8'hd5;
frames[14][1][25] = 8'hb1;
frames[14][1][26] = 8'h8d;
frames[14][1][27] = 8'h68;
frames[14][1][28] = 8'h24;
frames[14][1][29] = 8'h20;
frames[14][1][30] = 8'h00;
frames[14][1][31] = 8'h24;
frames[14][1][32] = 8'h24;
frames[14][1][33] = 8'h20;
frames[14][1][34] = 8'h24;
frames[14][1][35] = 8'h24;
frames[14][1][36] = 8'h91;
frames[14][1][37] = 8'hb6;
frames[14][1][38] = 8'hda;
frames[14][1][39] = 8'h6d;
frames[14][2][0] = 8'hd2;
frames[14][2][1] = 8'had;
frames[14][2][2] = 8'h89;
frames[14][2][3] = 8'had;
frames[14][2][4] = 8'h8d;
frames[14][2][5] = 8'h89;
frames[14][2][6] = 8'h89;
frames[14][2][7] = 8'h64;
frames[14][2][8] = 8'hb1;
frames[14][2][9] = 8'hfa;
frames[14][2][10] = 8'hd6;
frames[14][2][11] = 8'hd6;
frames[14][2][12] = 8'hd5;
frames[14][2][13] = 8'hd6;
frames[14][2][14] = 8'hd6;
frames[14][2][15] = 8'hd6;
frames[14][2][16] = 8'hd5;
frames[14][2][17] = 8'hd5;
frames[14][2][18] = 8'hd5;
frames[14][2][19] = 8'hd5;
frames[14][2][20] = 8'hd5;
frames[14][2][21] = 8'hd6;
frames[14][2][22] = 8'hd6;
frames[14][2][23] = 8'hb1;
frames[14][2][24] = 8'h69;
frames[14][2][25] = 8'h44;
frames[14][2][26] = 8'h24;
frames[14][2][27] = 8'h20;
frames[14][2][28] = 8'h24;
frames[14][2][29] = 8'h00;
frames[14][2][30] = 8'h00;
frames[14][2][31] = 8'h20;
frames[14][2][32] = 8'h20;
frames[14][2][33] = 8'h20;
frames[14][2][34] = 8'h20;
frames[14][2][35] = 8'h20;
frames[14][2][36] = 8'h6e;
frames[14][2][37] = 8'h6d;
frames[14][2][38] = 8'h4e;
frames[14][2][39] = 8'h72;
frames[14][3][0] = 8'hd6;
frames[14][3][1] = 8'had;
frames[14][3][2] = 8'h89;
frames[14][3][3] = 8'had;
frames[14][3][4] = 8'had;
frames[14][3][5] = 8'h88;
frames[14][3][6] = 8'h8d;
frames[14][3][7] = 8'h64;
frames[14][3][8] = 8'h8d;
frames[14][3][9] = 8'hb1;
frames[14][3][10] = 8'hd5;
frames[14][3][11] = 8'hd6;
frames[14][3][12] = 8'hd5;
frames[14][3][13] = 8'hd5;
frames[14][3][14] = 8'hd5;
frames[14][3][15] = 8'hd5;
frames[14][3][16] = 8'hd5;
frames[14][3][17] = 8'hb1;
frames[14][3][18] = 8'hd5;
frames[14][3][19] = 8'hd5;
frames[14][3][20] = 8'hb1;
frames[14][3][21] = 8'h8d;
frames[14][3][22] = 8'h69;
frames[14][3][23] = 8'h24;
frames[14][3][24] = 8'h20;
frames[14][3][25] = 8'h20;
frames[14][3][26] = 8'h24;
frames[14][3][27] = 8'h48;
frames[14][3][28] = 8'hb1;
frames[14][3][29] = 8'h8d;
frames[14][3][30] = 8'h48;
frames[14][3][31] = 8'h48;
frames[14][3][32] = 8'h69;
frames[14][3][33] = 8'h48;
frames[14][3][34] = 8'h48;
frames[14][3][35] = 8'h69;
frames[14][3][36] = 8'h8d;
frames[14][3][37] = 8'h69;
frames[14][3][38] = 8'h49;
frames[14][3][39] = 8'h6e;
frames[14][4][0] = 8'hf6;
frames[14][4][1] = 8'had;
frames[14][4][2] = 8'h89;
frames[14][4][3] = 8'had;
frames[14][4][4] = 8'had;
frames[14][4][5] = 8'h88;
frames[14][4][6] = 8'h88;
frames[14][4][7] = 8'h88;
frames[14][4][8] = 8'h64;
frames[14][4][9] = 8'h64;
frames[14][4][10] = 8'h68;
frames[14][4][11] = 8'hd1;
frames[14][4][12] = 8'hd1;
frames[14][4][13] = 8'hd1;
frames[14][4][14] = 8'hb1;
frames[14][4][15] = 8'hd5;
frames[14][4][16] = 8'hb6;
frames[14][4][17] = 8'hb1;
frames[14][4][18] = 8'h91;
frames[14][4][19] = 8'h6d;
frames[14][4][20] = 8'h44;
frames[14][4][21] = 8'h24;
frames[14][4][22] = 8'h24;
frames[14][4][23] = 8'h20;
frames[14][4][24] = 8'h44;
frames[14][4][25] = 8'h6d;
frames[14][4][26] = 8'hb1;
frames[14][4][27] = 8'hb6;
frames[14][4][28] = 8'hd6;
frames[14][4][29] = 8'hd6;
frames[14][4][30] = 8'hb6;
frames[14][4][31] = 8'hb5;
frames[14][4][32] = 8'hb5;
frames[14][4][33] = 8'hb1;
frames[14][4][34] = 8'hb1;
frames[14][4][35] = 8'hb1;
frames[14][4][36] = 8'hb6;
frames[14][4][37] = 8'h8d;
frames[14][4][38] = 8'h8d;
frames[14][4][39] = 8'h6d;
frames[14][5][0] = 8'hf6;
frames[14][5][1] = 8'had;
frames[14][5][2] = 8'ha9;
frames[14][5][3] = 8'h89;
frames[14][5][4] = 8'had;
frames[14][5][5] = 8'h89;
frames[14][5][6] = 8'h64;
frames[14][5][7] = 8'h88;
frames[14][5][8] = 8'h88;
frames[14][5][9] = 8'h89;
frames[14][5][10] = 8'had;
frames[14][5][11] = 8'hd1;
frames[14][5][12] = 8'hb2;
frames[14][5][13] = 8'hb1;
frames[14][5][14] = 8'hb2;
frames[14][5][15] = 8'hb1;
frames[14][5][16] = 8'h8d;
frames[14][5][17] = 8'h48;
frames[14][5][18] = 8'h24;
frames[14][5][19] = 8'h24;
frames[14][5][20] = 8'h24;
frames[14][5][21] = 8'h24;
frames[14][5][22] = 8'h24;
frames[14][5][23] = 8'h49;
frames[14][5][24] = 8'hb1;
frames[14][5][25] = 8'hd6;
frames[14][5][26] = 8'hd5;
frames[14][5][27] = 8'hd6;
frames[14][5][28] = 8'hd5;
frames[14][5][29] = 8'hd5;
frames[14][5][30] = 8'hb5;
frames[14][5][31] = 8'hb5;
frames[14][5][32] = 8'hd6;
frames[14][5][33] = 8'hb5;
frames[14][5][34] = 8'hb1;
frames[14][5][35] = 8'hb1;
frames[14][5][36] = 8'hb1;
frames[14][5][37] = 8'hd6;
frames[14][5][38] = 8'hb6;
frames[14][5][39] = 8'h6d;
frames[14][6][0] = 8'hfb;
frames[14][6][1] = 8'hb1;
frames[14][6][2] = 8'had;
frames[14][6][3] = 8'h88;
frames[14][6][4] = 8'h88;
frames[14][6][5] = 8'had;
frames[14][6][6] = 8'h89;
frames[14][6][7] = 8'h64;
frames[14][6][8] = 8'h8d;
frames[14][6][9] = 8'had;
frames[14][6][10] = 8'hd6;
frames[14][6][11] = 8'hd6;
frames[14][6][12] = 8'hd6;
frames[14][6][13] = 8'hb1;
frames[14][6][14] = 8'h69;
frames[14][6][15] = 8'h24;
frames[14][6][16] = 8'h24;
frames[14][6][17] = 8'h24;
frames[14][6][18] = 8'h24;
frames[14][6][19] = 8'h24;
frames[14][6][20] = 8'h24;
frames[14][6][21] = 8'h44;
frames[14][6][22] = 8'h8d;
frames[14][6][23] = 8'hb6;
frames[14][6][24] = 8'hb1;
frames[14][6][25] = 8'hb1;
frames[14][6][26] = 8'hb1;
frames[14][6][27] = 8'hb5;
frames[14][6][28] = 8'hd5;
frames[14][6][29] = 8'hd5;
frames[14][6][30] = 8'hd5;
frames[14][6][31] = 8'hd5;
frames[14][6][32] = 8'hb5;
frames[14][6][33] = 8'hb1;
frames[14][6][34] = 8'hb1;
frames[14][6][35] = 8'h91;
frames[14][6][36] = 8'h8d;
frames[14][6][37] = 8'hb1;
frames[14][6][38] = 8'h8d;
frames[14][6][39] = 8'h68;
frames[14][7][0] = 8'hff;
frames[14][7][1] = 8'hfa;
frames[14][7][2] = 8'hb1;
frames[14][7][3] = 8'had;
frames[14][7][4] = 8'h88;
frames[14][7][5] = 8'had;
frames[14][7][6] = 8'had;
frames[14][7][7] = 8'h88;
frames[14][7][8] = 8'h64;
frames[14][7][9] = 8'h88;
frames[14][7][10] = 8'hb2;
frames[14][7][11] = 8'h8d;
frames[14][7][12] = 8'h48;
frames[14][7][13] = 8'h24;
frames[14][7][14] = 8'h24;
frames[14][7][15] = 8'h24;
frames[14][7][16] = 8'h24;
frames[14][7][17] = 8'h20;
frames[14][7][18] = 8'h20;
frames[14][7][19] = 8'h24;
frames[14][7][20] = 8'h6d;
frames[14][7][21] = 8'hb6;
frames[14][7][22] = 8'hd6;
frames[14][7][23] = 8'hd6;
frames[14][7][24] = 8'hb1;
frames[14][7][25] = 8'hd6;
frames[14][7][26] = 8'hb5;
frames[14][7][27] = 8'hb5;
frames[14][7][28] = 8'hd5;
frames[14][7][29] = 8'hd6;
frames[14][7][30] = 8'hd6;
frames[14][7][31] = 8'hd6;
frames[14][7][32] = 8'hd6;
frames[14][7][33] = 8'hb5;
frames[14][7][34] = 8'hb1;
frames[14][7][35] = 8'hb1;
frames[14][7][36] = 8'h91;
frames[14][7][37] = 8'hb1;
frames[14][7][38] = 8'hb1;
frames[14][7][39] = 8'h8d;
frames[14][8][0] = 8'hfa;
frames[14][8][1] = 8'hff;
frames[14][8][2] = 8'hf6;
frames[14][8][3] = 8'had;
frames[14][8][4] = 8'had;
frames[14][8][5] = 8'had;
frames[14][8][6] = 8'had;
frames[14][8][7] = 8'had;
frames[14][8][8] = 8'h88;
frames[14][8][9] = 8'h88;
frames[14][8][10] = 8'h68;
frames[14][8][11] = 8'h44;
frames[14][8][12] = 8'h24;
frames[14][8][13] = 8'h24;
frames[14][8][14] = 8'h24;
frames[14][8][15] = 8'h24;
frames[14][8][16] = 8'h24;
frames[14][8][17] = 8'h48;
frames[14][8][18] = 8'h6d;
frames[14][8][19] = 8'hb2;
frames[14][8][20] = 8'hd6;
frames[14][8][21] = 8'hd6;
frames[14][8][22] = 8'hd6;
frames[14][8][23] = 8'hd6;
frames[14][8][24] = 8'hd5;
frames[14][8][25] = 8'hd5;
frames[14][8][26] = 8'hd5;
frames[14][8][27] = 8'hd5;
frames[14][8][28] = 8'hd6;
frames[14][8][29] = 8'hd6;
frames[14][8][30] = 8'hd6;
frames[14][8][31] = 8'hb5;
frames[14][8][32] = 8'hb5;
frames[14][8][33] = 8'hb1;
frames[14][8][34] = 8'hb1;
frames[14][8][35] = 8'hb1;
frames[14][8][36] = 8'hb5;
frames[14][8][37] = 8'hb1;
frames[14][8][38] = 8'hb2;
frames[14][8][39] = 8'h91;
frames[14][9][0] = 8'hff;
frames[14][9][1] = 8'hff;
frames[14][9][2] = 8'hff;
frames[14][9][3] = 8'hb2;
frames[14][9][4] = 8'ha9;
frames[14][9][5] = 8'h89;
frames[14][9][6] = 8'h88;
frames[14][9][7] = 8'had;
frames[14][9][8] = 8'hb1;
frames[14][9][9] = 8'hb1;
frames[14][9][10] = 8'h8d;
frames[14][9][11] = 8'h68;
frames[14][9][12] = 8'h48;
frames[14][9][13] = 8'h44;
frames[14][9][14] = 8'h48;
frames[14][9][15] = 8'h6d;
frames[14][9][16] = 8'h91;
frames[14][9][17] = 8'hb6;
frames[14][9][18] = 8'hb6;
frames[14][9][19] = 8'hb6;
frames[14][9][20] = 8'hd5;
frames[14][9][21] = 8'hd5;
frames[14][9][22] = 8'hd6;
frames[14][9][23] = 8'hd5;
frames[14][9][24] = 8'hd5;
frames[14][9][25] = 8'hb1;
frames[14][9][26] = 8'hb1;
frames[14][9][27] = 8'hb1;
frames[14][9][28] = 8'hb5;
frames[14][9][29] = 8'hd5;
frames[14][9][30] = 8'hb5;
frames[14][9][31] = 8'hb1;
frames[14][9][32] = 8'h8d;
frames[14][9][33] = 8'h68;
frames[14][9][34] = 8'h68;
frames[14][9][35] = 8'had;
frames[14][9][36] = 8'hb1;
frames[14][9][37] = 8'hb1;
frames[14][9][38] = 8'hb1;
frames[14][9][39] = 8'h8d;
frames[14][10][0] = 8'hff;
frames[14][10][1] = 8'hfb;
frames[14][10][2] = 8'hb6;
frames[14][10][3] = 8'h6d;
frames[14][10][4] = 8'h88;
frames[14][10][5] = 8'had;
frames[14][10][6] = 8'h88;
frames[14][10][7] = 8'had;
frames[14][10][8] = 8'hb1;
frames[14][10][9] = 8'hd5;
frames[14][10][10] = 8'hb1;
frames[14][10][11] = 8'h8d;
frames[14][10][12] = 8'h8d;
frames[14][10][13] = 8'hb2;
frames[14][10][14] = 8'hb6;
frames[14][10][15] = 8'hd6;
frames[14][10][16] = 8'hd6;
frames[14][10][17] = 8'hb6;
frames[14][10][18] = 8'hb5;
frames[14][10][19] = 8'hb5;
frames[14][10][20] = 8'hd5;
frames[14][10][21] = 8'hd5;
frames[14][10][22] = 8'hd5;
frames[14][10][23] = 8'hb1;
frames[14][10][24] = 8'hd6;
frames[14][10][25] = 8'had;
frames[14][10][26] = 8'h8d;
frames[14][10][27] = 8'h8d;
frames[14][10][28] = 8'hb1;
frames[14][10][29] = 8'h91;
frames[14][10][30] = 8'h91;
frames[14][10][31] = 8'hb1;
frames[14][10][32] = 8'h91;
frames[14][10][33] = 8'h91;
frames[14][10][34] = 8'h8d;
frames[14][10][35] = 8'hb1;
frames[14][10][36] = 8'hd6;
frames[14][10][37] = 8'h8d;
frames[14][10][38] = 8'h68;
frames[14][10][39] = 8'h48;
frames[14][11][0] = 8'h6d;
frames[14][11][1] = 8'h44;
frames[14][11][2] = 8'h24;
frames[14][11][3] = 8'h24;
frames[14][11][4] = 8'h69;
frames[14][11][5] = 8'hb6;
frames[14][11][6] = 8'hb1;
frames[14][11][7] = 8'hd1;
frames[14][11][8] = 8'hd1;
frames[14][11][9] = 8'hb1;
frames[14][11][10] = 8'hb1;
frames[14][11][11] = 8'hb1;
frames[14][11][12] = 8'hb6;
frames[14][11][13] = 8'hb6;
frames[14][11][14] = 8'hb6;
frames[14][11][15] = 8'hd6;
frames[14][11][16] = 8'hd6;
frames[14][11][17] = 8'hd6;
frames[14][11][18] = 8'hb2;
frames[14][11][19] = 8'h8d;
frames[14][11][20] = 8'hb1;
frames[14][11][21] = 8'hb1;
frames[14][11][22] = 8'hd5;
frames[14][11][23] = 8'hd5;
frames[14][11][24] = 8'hb1;
frames[14][11][25] = 8'h8d;
frames[14][11][26] = 8'h8d;
frames[14][11][27] = 8'h8d;
frames[14][11][28] = 8'hb1;
frames[14][11][29] = 8'hb1;
frames[14][11][30] = 8'hb1;
frames[14][11][31] = 8'hb1;
frames[14][11][32] = 8'hb1;
frames[14][11][33] = 8'h91;
frames[14][11][34] = 8'h8d;
frames[14][11][35] = 8'h8d;
frames[14][11][36] = 8'hb1;
frames[14][11][37] = 8'h48;
frames[14][11][38] = 8'h44;
frames[14][11][39] = 8'h44;
frames[14][12][0] = 8'h24;
frames[14][12][1] = 8'h24;
frames[14][12][2] = 8'h44;
frames[14][12][3] = 8'h44;
frames[14][12][4] = 8'h68;
frames[14][12][5] = 8'hd6;
frames[14][12][6] = 8'hb1;
frames[14][12][7] = 8'hb1;
frames[14][12][8] = 8'hb1;
frames[14][12][9] = 8'hd1;
frames[14][12][10] = 8'hd5;
frames[14][12][11] = 8'hb1;
frames[14][12][12] = 8'hb1;
frames[14][12][13] = 8'hb1;
frames[14][12][14] = 8'hb1;
frames[14][12][15] = 8'h88;
frames[14][12][16] = 8'h8d;
frames[14][12][17] = 8'hd2;
frames[14][12][18] = 8'h91;
frames[14][12][19] = 8'h44;
frames[14][12][20] = 8'h24;
frames[14][12][21] = 8'h48;
frames[14][12][22] = 8'h8d;
frames[14][12][23] = 8'h91;
frames[14][12][24] = 8'h8d;
frames[14][12][25] = 8'h8d;
frames[14][12][26] = 8'h69;
frames[14][12][27] = 8'h69;
frames[14][12][28] = 8'h8d;
frames[14][12][29] = 8'h8d;
frames[14][12][30] = 8'h69;
frames[14][12][31] = 8'h68;
frames[14][12][32] = 8'h48;
frames[14][12][33] = 8'h48;
frames[14][12][34] = 8'h44;
frames[14][12][35] = 8'h69;
frames[14][12][36] = 8'hb2;
frames[14][12][37] = 8'h69;
frames[14][12][38] = 8'h44;
frames[14][12][39] = 8'h44;
frames[14][13][0] = 8'h68;
frames[14][13][1] = 8'h69;
frames[14][13][2] = 8'had;
frames[14][13][3] = 8'hd1;
frames[14][13][4] = 8'had;
frames[14][13][5] = 8'hd1;
frames[14][13][6] = 8'h8d;
frames[14][13][7] = 8'had;
frames[14][13][8] = 8'hb1;
frames[14][13][9] = 8'hb1;
frames[14][13][10] = 8'hb1;
frames[14][13][11] = 8'hb1;
frames[14][13][12] = 8'hb1;
frames[14][13][13] = 8'hb1;
frames[14][13][14] = 8'hd1;
frames[14][13][15] = 8'hb1;
frames[14][13][16] = 8'h64;
frames[14][13][17] = 8'h88;
frames[14][13][18] = 8'hb2;
frames[14][13][19] = 8'h8d;
frames[14][13][20] = 8'h44;
frames[14][13][21] = 8'h24;
frames[14][13][22] = 8'h8d;
frames[14][13][23] = 8'h8d;
frames[14][13][24] = 8'h69;
frames[14][13][25] = 8'h6d;
frames[14][13][26] = 8'h8d;
frames[14][13][27] = 8'h6d;
frames[14][13][28] = 8'h6d;
frames[14][13][29] = 8'h6d;
frames[14][13][30] = 8'h6d;
frames[14][13][31] = 8'h6d;
frames[14][13][32] = 8'h6d;
frames[14][13][33] = 8'h6d;
frames[14][13][34] = 8'h6d;
frames[14][13][35] = 8'h8d;
frames[14][13][36] = 8'hb6;
frames[14][13][37] = 8'h8d;
frames[14][13][38] = 8'h68;
frames[14][13][39] = 8'h48;
frames[14][14][0] = 8'hd6;
frames[14][14][1] = 8'hd6;
frames[14][14][2] = 8'hd1;
frames[14][14][3] = 8'had;
frames[14][14][4] = 8'hb1;
frames[14][14][5] = 8'hd5;
frames[14][14][6] = 8'had;
frames[14][14][7] = 8'h8d;
frames[14][14][8] = 8'h8d;
frames[14][14][9] = 8'hd5;
frames[14][14][10] = 8'hb5;
frames[14][14][11] = 8'hb5;
frames[14][14][12] = 8'hb1;
frames[14][14][13] = 8'hb1;
frames[14][14][14] = 8'hb1;
frames[14][14][15] = 8'hb1;
frames[14][14][16] = 8'hb1;
frames[14][14][17] = 8'h88;
frames[14][14][18] = 8'hb1;
frames[14][14][19] = 8'hd6;
frames[14][14][20] = 8'hb2;
frames[14][14][21] = 8'h8d;
frames[14][14][22] = 8'hb6;
frames[14][14][23] = 8'hb6;
frames[14][14][24] = 8'hb2;
frames[14][14][25] = 8'hb2;
frames[14][14][26] = 8'hb2;
frames[14][14][27] = 8'h91;
frames[14][14][28] = 8'h8d;
frames[14][14][29] = 8'h8d;
frames[14][14][30] = 8'h8d;
frames[14][14][31] = 8'h8d;
frames[14][14][32] = 8'h8d;
frames[14][14][33] = 8'h6d;
frames[14][14][34] = 8'h6d;
frames[14][14][35] = 8'h6d;
frames[14][14][36] = 8'hb2;
frames[14][14][37] = 8'h91;
frames[14][14][38] = 8'h6d;
frames[14][14][39] = 8'h6d;
frames[14][15][0] = 8'hd6;
frames[14][15][1] = 8'hd6;
frames[14][15][2] = 8'hb1;
frames[14][15][3] = 8'hb1;
frames[14][15][4] = 8'hb1;
frames[14][15][5] = 8'hb1;
frames[14][15][6] = 8'hb1;
frames[14][15][7] = 8'h8c;
frames[14][15][8] = 8'hd5;
frames[14][15][9] = 8'hd6;
frames[14][15][10] = 8'hd5;
frames[14][15][11] = 8'hb5;
frames[14][15][12] = 8'hb1;
frames[14][15][13] = 8'h8d;
frames[14][15][14] = 8'h8d;
frames[14][15][15] = 8'h68;
frames[14][15][16] = 8'h8d;
frames[14][15][17] = 8'had;
frames[14][15][18] = 8'hb1;
frames[14][15][19] = 8'hb1;
frames[14][15][20] = 8'hb1;
frames[14][15][21] = 8'h8d;
frames[14][15][22] = 8'hb6;
frames[14][15][23] = 8'hb6;
frames[14][15][24] = 8'hb2;
frames[14][15][25] = 8'h91;
frames[14][15][26] = 8'h8d;
frames[14][15][27] = 8'h91;
frames[14][15][28] = 8'h8d;
frames[14][15][29] = 8'h8d;
frames[14][15][30] = 8'h8d;
frames[14][15][31] = 8'h8d;
frames[14][15][32] = 8'h69;
frames[14][15][33] = 8'h44;
frames[14][15][34] = 8'h24;
frames[14][15][35] = 8'h6d;
frames[14][15][36] = 8'hff;
frames[14][15][37] = 8'h91;
frames[14][15][38] = 8'h44;
frames[14][15][39] = 8'h44;
frames[14][16][0] = 8'hd5;
frames[14][16][1] = 8'hd5;
frames[14][16][2] = 8'hd6;
frames[14][16][3] = 8'hd6;
frames[14][16][4] = 8'hb1;
frames[14][16][5] = 8'h8c;
frames[14][16][6] = 8'hb1;
frames[14][16][7] = 8'had;
frames[14][16][8] = 8'hb1;
frames[14][16][9] = 8'hb1;
frames[14][16][10] = 8'hb1;
frames[14][16][11] = 8'h8d;
frames[14][16][12] = 8'hb1;
frames[14][16][13] = 8'hb1;
frames[14][16][14] = 8'hb1;
frames[14][16][15] = 8'h68;
frames[14][16][16] = 8'h64;
frames[14][16][17] = 8'had;
frames[14][16][18] = 8'h8d;
frames[14][16][19] = 8'hb1;
frames[14][16][20] = 8'hb1;
frames[14][16][21] = 8'hb1;
frames[14][16][22] = 8'hb2;
frames[14][16][23] = 8'hb2;
frames[14][16][24] = 8'h91;
frames[14][16][25] = 8'hb2;
frames[14][16][26] = 8'hb6;
frames[14][16][27] = 8'hb6;
frames[14][16][28] = 8'h92;
frames[14][16][29] = 8'h91;
frames[14][16][30] = 8'h6d;
frames[14][16][31] = 8'h48;
frames[14][16][32] = 8'h24;
frames[14][16][33] = 8'h24;
frames[14][16][34] = 8'h24;
frames[14][16][35] = 8'h69;
frames[14][16][36] = 8'hb6;
frames[14][16][37] = 8'h6d;
frames[14][16][38] = 8'h44;
frames[14][16][39] = 8'h44;
frames[14][17][0] = 8'hd5;
frames[14][17][1] = 8'hb1;
frames[14][17][2] = 8'hb1;
frames[14][17][3] = 8'had;
frames[14][17][4] = 8'h8d;
frames[14][17][5] = 8'h68;
frames[14][17][6] = 8'h8d;
frames[14][17][7] = 8'hd6;
frames[14][17][8] = 8'h8d;
frames[14][17][9] = 8'h88;
frames[14][17][10] = 8'hb1;
frames[14][17][11] = 8'h8d;
frames[14][17][12] = 8'h8d;
frames[14][17][13] = 8'hb1;
frames[14][17][14] = 8'had;
frames[14][17][15] = 8'h8d;
frames[14][17][16] = 8'h64;
frames[14][17][17] = 8'h89;
frames[14][17][18] = 8'h8d;
frames[14][17][19] = 8'hd6;
frames[14][17][20] = 8'h8d;
frames[14][17][21] = 8'h91;
frames[14][17][22] = 8'hb2;
frames[14][17][23] = 8'hb6;
frames[14][17][24] = 8'hb6;
frames[14][17][25] = 8'hb6;
frames[14][17][26] = 8'hd6;
frames[14][17][27] = 8'hb6;
frames[14][17][28] = 8'h6d;
frames[14][17][29] = 8'h49;
frames[14][17][30] = 8'h24;
frames[14][17][31] = 8'h24;
frames[14][17][32] = 8'h24;
frames[14][17][33] = 8'h24;
frames[14][17][34] = 8'h44;
frames[14][17][35] = 8'h48;
frames[14][17][36] = 8'h44;
frames[14][17][37] = 8'h44;
frames[14][17][38] = 8'h44;
frames[14][17][39] = 8'h44;
frames[14][18][0] = 8'had;
frames[14][18][1] = 8'h88;
frames[14][18][2] = 8'h88;
frames[14][18][3] = 8'had;
frames[14][18][4] = 8'hd5;
frames[14][18][5] = 8'hd5;
frames[14][18][6] = 8'hb1;
frames[14][18][7] = 8'hd1;
frames[14][18][8] = 8'ha8;
frames[14][18][9] = 8'h84;
frames[14][18][10] = 8'h88;
frames[14][18][11] = 8'had;
frames[14][18][12] = 8'hb5;
frames[14][18][13] = 8'hb1;
frames[14][18][14] = 8'h8d;
frames[14][18][15] = 8'hb1;
frames[14][18][16] = 8'h8d;
frames[14][18][17] = 8'h68;
frames[14][18][18] = 8'h8d;
frames[14][18][19] = 8'h8d;
frames[14][18][20] = 8'h69;
frames[14][18][21] = 8'h6d;
frames[14][18][22] = 8'h91;
frames[14][18][23] = 8'hb6;
frames[14][18][24] = 8'hb6;
frames[14][18][25] = 8'hb2;
frames[14][18][26] = 8'h8d;
frames[14][18][27] = 8'h6d;
frames[14][18][28] = 8'h44;
frames[14][18][29] = 8'h24;
frames[14][18][30] = 8'h24;
frames[14][18][31] = 8'h24;
frames[14][18][32] = 8'h44;
frames[14][18][33] = 8'h44;
frames[14][18][34] = 8'h48;
frames[14][18][35] = 8'h69;
frames[14][18][36] = 8'h6d;
frames[14][18][37] = 8'h68;
frames[14][18][38] = 8'h68;
frames[14][18][39] = 8'h8d;
frames[14][19][0] = 8'hb1;
frames[14][19][1] = 8'hb1;
frames[14][19][2] = 8'hb1;
frames[14][19][3] = 8'hd6;
frames[14][19][4] = 8'hb1;
frames[14][19][5] = 8'hd6;
frames[14][19][6] = 8'hd6;
frames[14][19][7] = 8'hb1;
frames[14][19][8] = 8'hb1;
frames[14][19][9] = 8'h8d;
frames[14][19][10] = 8'h88;
frames[14][19][11] = 8'h88;
frames[14][19][12] = 8'hb1;
frames[14][19][13] = 8'hb5;
frames[14][19][14] = 8'hb1;
frames[14][19][15] = 8'hb1;
frames[14][19][16] = 8'hb1;
frames[14][19][17] = 8'h8d;
frames[14][19][18] = 8'h69;
frames[14][19][19] = 8'h91;
frames[14][19][20] = 8'hb6;
frames[14][19][21] = 8'h69;
frames[14][19][22] = 8'h69;
frames[14][19][23] = 8'h8d;
frames[14][19][24] = 8'h91;
frames[14][19][25] = 8'h8d;
frames[14][19][26] = 8'h8d;
frames[14][19][27] = 8'h6d;
frames[14][19][28] = 8'h6d;
frames[14][19][29] = 8'h6d;
frames[14][19][30] = 8'h68;
frames[14][19][31] = 8'h68;
frames[14][19][32] = 8'h68;
frames[14][19][33] = 8'h68;
frames[14][19][34] = 8'h8d;
frames[14][19][35] = 8'h8d;
frames[14][19][36] = 8'h8d;
frames[14][19][37] = 8'h8d;
frames[14][19][38] = 8'h8d;
frames[14][19][39] = 8'h8d;
frames[14][20][0] = 8'hb1;
frames[14][20][1] = 8'h91;
frames[14][20][2] = 8'hb1;
frames[14][20][3] = 8'hb1;
frames[14][20][4] = 8'hb1;
frames[14][20][5] = 8'hb5;
frames[14][20][6] = 8'hb6;
frames[14][20][7] = 8'hd6;
frames[14][20][8] = 8'hd6;
frames[14][20][9] = 8'hb1;
frames[14][20][10] = 8'hb5;
frames[14][20][11] = 8'hb1;
frames[14][20][12] = 8'hb1;
frames[14][20][13] = 8'hb1;
frames[14][20][14] = 8'hb6;
frames[14][20][15] = 8'h8d;
frames[14][20][16] = 8'h48;
frames[14][20][17] = 8'h6d;
frames[14][20][18] = 8'hb6;
frames[14][20][19] = 8'hd6;
frames[14][20][20] = 8'hb2;
frames[14][20][21] = 8'h69;
frames[14][20][22] = 8'h68;
frames[14][20][23] = 8'h68;
frames[14][20][24] = 8'h68;
frames[14][20][25] = 8'h69;
frames[14][20][26] = 8'h68;
frames[14][20][27] = 8'h8d;
frames[14][20][28] = 8'h8d;
frames[14][20][29] = 8'hb6;
frames[14][20][30] = 8'hb1;
frames[14][20][31] = 8'h8d;
frames[14][20][32] = 8'had;
frames[14][20][33] = 8'had;
frames[14][20][34] = 8'had;
frames[14][20][35] = 8'hb1;
frames[14][20][36] = 8'hb1;
frames[14][20][37] = 8'hb1;
frames[14][20][38] = 8'hb1;
frames[14][20][39] = 8'hb1;
frames[14][21][0] = 8'h44;
frames[14][21][1] = 8'h68;
frames[14][21][2] = 8'h6d;
frames[14][21][3] = 8'h8d;
frames[14][21][4] = 8'h91;
frames[14][21][5] = 8'hb1;
frames[14][21][6] = 8'hb1;
frames[14][21][7] = 8'hb1;
frames[14][21][8] = 8'hb1;
frames[14][21][9] = 8'hb1;
frames[14][21][10] = 8'h8d;
frames[14][21][11] = 8'h8d;
frames[14][21][12] = 8'h6d;
frames[14][21][13] = 8'h6d;
frames[14][21][14] = 8'h91;
frames[14][21][15] = 8'h8d;
frames[14][21][16] = 8'hb2;
frames[14][21][17] = 8'hd6;
frames[14][21][18] = 8'h92;
frames[14][21][19] = 8'h49;
frames[14][21][20] = 8'h44;
frames[14][21][21] = 8'h48;
frames[14][21][22] = 8'h69;
frames[14][21][23] = 8'h69;
frames[14][21][24] = 8'h8d;
frames[14][21][25] = 8'hb1;
frames[14][21][26] = 8'hb1;
frames[14][21][27] = 8'hb1;
frames[14][21][28] = 8'hb1;
frames[14][21][29] = 8'hd6;
frames[14][21][30] = 8'hd6;
frames[14][21][31] = 8'hd6;
frames[14][21][32] = 8'hd6;
frames[14][21][33] = 8'hd6;
frames[14][21][34] = 8'hd5;
frames[14][21][35] = 8'hd6;
frames[14][21][36] = 8'hd5;
frames[14][21][37] = 8'hd5;
frames[14][21][38] = 8'hb5;
frames[14][21][39] = 8'hb1;
frames[14][22][0] = 8'hb2;
frames[14][22][1] = 8'h49;
frames[14][22][2] = 8'h20;
frames[14][22][3] = 8'h20;
frames[14][22][4] = 8'h24;
frames[14][22][5] = 8'h24;
frames[14][22][6] = 8'h24;
frames[14][22][7] = 8'h24;
frames[14][22][8] = 8'h24;
frames[14][22][9] = 8'h24;
frames[14][22][10] = 8'h24;
frames[14][22][11] = 8'h44;
frames[14][22][12] = 8'h6d;
frames[14][22][13] = 8'hb6;
frames[14][22][14] = 8'hd6;
frames[14][22][15] = 8'hb6;
frames[14][22][16] = 8'h8d;
frames[14][22][17] = 8'h48;
frames[14][22][18] = 8'h24;
frames[14][22][19] = 8'h20;
frames[14][22][20] = 8'h20;
frames[14][22][21] = 8'h44;
frames[14][22][22] = 8'h68;
frames[14][22][23] = 8'h8d;
frames[14][22][24] = 8'h91;
frames[14][22][25] = 8'hd6;
frames[14][22][26] = 8'hda;
frames[14][22][27] = 8'hb6;
frames[14][22][28] = 8'hb6;
frames[14][22][29] = 8'hd6;
frames[14][22][30] = 8'hd6;
frames[14][22][31] = 8'hd6;
frames[14][22][32] = 8'hd5;
frames[14][22][33] = 8'hd5;
frames[14][22][34] = 8'hd5;
frames[14][22][35] = 8'hd5;
frames[14][22][36] = 8'hb5;
frames[14][22][37] = 8'hb1;
frames[14][22][38] = 8'hb1;
frames[14][22][39] = 8'hb1;
frames[14][23][0] = 8'hb2;
frames[14][23][1] = 8'hb6;
frames[14][23][2] = 8'h6d;
frames[14][23][3] = 8'h44;
frames[14][23][4] = 8'h24;
frames[14][23][5] = 8'h24;
frames[14][23][6] = 8'h24;
frames[14][23][7] = 8'h24;
frames[14][23][8] = 8'h24;
frames[14][23][9] = 8'h44;
frames[14][23][10] = 8'h6d;
frames[14][23][11] = 8'h8d;
frames[14][23][12] = 8'hb2;
frames[14][23][13] = 8'h92;
frames[14][23][14] = 8'h6d;
frames[14][23][15] = 8'h24;
frames[14][23][16] = 8'h24;
frames[14][23][17] = 8'h20;
frames[14][23][18] = 8'h20;
frames[14][23][19] = 8'h24;
frames[14][23][20] = 8'h20;
frames[14][23][21] = 8'h44;
frames[14][23][22] = 8'h68;
frames[14][23][23] = 8'h8d;
frames[14][23][24] = 8'h8d;
frames[14][23][25] = 8'h8d;
frames[14][23][26] = 8'hb1;
frames[14][23][27] = 8'hb1;
frames[14][23][28] = 8'hb1;
frames[14][23][29] = 8'hb1;
frames[14][23][30] = 8'hb1;
frames[14][23][31] = 8'hb1;
frames[14][23][32] = 8'hb1;
frames[14][23][33] = 8'hb1;
frames[14][23][34] = 8'hb1;
frames[14][23][35] = 8'hb1;
frames[14][23][36] = 8'hb1;
frames[14][23][37] = 8'hb1;
frames[14][23][38] = 8'hb1;
frames[14][23][39] = 8'hb5;
frames[14][24][0] = 8'h44;
frames[14][24][1] = 8'h44;
frames[14][24][2] = 8'h69;
frames[14][24][3] = 8'h69;
frames[14][24][4] = 8'h44;
frames[14][24][5] = 8'h44;
frames[14][24][6] = 8'h44;
frames[14][24][7] = 8'h44;
frames[14][24][8] = 8'h44;
frames[14][24][9] = 8'h49;
frames[14][24][10] = 8'h69;
frames[14][24][11] = 8'h69;
frames[14][24][12] = 8'h44;
frames[14][24][13] = 8'h24;
frames[14][24][14] = 8'h20;
frames[14][24][15] = 8'h20;
frames[14][24][16] = 8'h20;
frames[14][24][17] = 8'h20;
frames[14][24][18] = 8'h24;
frames[14][24][19] = 8'h44;
frames[14][24][20] = 8'h44;
frames[14][24][21] = 8'h44;
frames[14][24][22] = 8'h68;
frames[14][24][23] = 8'h8d;
frames[14][24][24] = 8'hd6;
frames[14][24][25] = 8'hd6;
frames[14][24][26] = 8'hb5;
frames[14][24][27] = 8'hb5;
frames[14][24][28] = 8'hb5;
frames[14][24][29] = 8'hb5;
frames[14][24][30] = 8'hb5;
frames[14][24][31] = 8'hb1;
frames[14][24][32] = 8'hb1;
frames[14][24][33] = 8'hb1;
frames[14][24][34] = 8'hb1;
frames[14][24][35] = 8'hd5;
frames[14][24][36] = 8'hd5;
frames[14][24][37] = 8'hd5;
frames[14][24][38] = 8'hd6;
frames[14][24][39] = 8'hd6;
frames[14][25][0] = 8'h44;
frames[14][25][1] = 8'h44;
frames[14][25][2] = 8'h24;
frames[14][25][3] = 8'h44;
frames[14][25][4] = 8'h44;
frames[14][25][5] = 8'h44;
frames[14][25][6] = 8'h44;
frames[14][25][7] = 8'h44;
frames[14][25][8] = 8'h44;
frames[14][25][9] = 8'h24;
frames[14][25][10] = 8'h24;
frames[14][25][11] = 8'h24;
frames[14][25][12] = 8'h20;
frames[14][25][13] = 8'h20;
frames[14][25][14] = 8'h20;
frames[14][25][15] = 8'h20;
frames[14][25][16] = 8'h24;
frames[14][25][17] = 8'h24;
frames[14][25][18] = 8'h44;
frames[14][25][19] = 8'h44;
frames[14][25][20] = 8'h64;
frames[14][25][21] = 8'h68;
frames[14][25][22] = 8'h88;
frames[14][25][23] = 8'had;
frames[14][25][24] = 8'hd6;
frames[14][25][25] = 8'hff;
frames[14][25][26] = 8'hda;
frames[14][25][27] = 8'hb5;
frames[14][25][28] = 8'hb5;
frames[14][25][29] = 8'hd5;
frames[14][25][30] = 8'hd5;
frames[14][25][31] = 8'hb5;
frames[14][25][32] = 8'hb5;
frames[14][25][33] = 8'hd5;
frames[14][25][34] = 8'hb5;
frames[14][25][35] = 8'hd5;
frames[14][25][36] = 8'hd5;
frames[14][25][37] = 8'hd5;
frames[14][25][38] = 8'hd6;
frames[14][25][39] = 8'hd6;
frames[14][26][0] = 8'h44;
frames[14][26][1] = 8'h24;
frames[14][26][2] = 8'h24;
frames[14][26][3] = 8'h24;
frames[14][26][4] = 8'h24;
frames[14][26][5] = 8'h24;
frames[14][26][6] = 8'h24;
frames[14][26][7] = 8'h44;
frames[14][26][8] = 8'h24;
frames[14][26][9] = 8'h24;
frames[14][26][10] = 8'h20;
frames[14][26][11] = 8'h24;
frames[14][26][12] = 8'h20;
frames[14][26][13] = 8'h24;
frames[14][26][14] = 8'h44;
frames[14][26][15] = 8'h44;
frames[14][26][16] = 8'h44;
frames[14][26][17] = 8'h44;
frames[14][26][18] = 8'h68;
frames[14][26][19] = 8'h68;
frames[14][26][20] = 8'h68;
frames[14][26][21] = 8'h8d;
frames[14][26][22] = 8'had;
frames[14][26][23] = 8'hb1;
frames[14][26][24] = 8'hb1;
frames[14][26][25] = 8'hd6;
frames[14][26][26] = 8'hd6;
frames[14][26][27] = 8'hb5;
frames[14][26][28] = 8'hd5;
frames[14][26][29] = 8'hb1;
frames[14][26][30] = 8'hb5;
frames[14][26][31] = 8'hb5;
frames[14][26][32] = 8'hb5;
frames[14][26][33] = 8'hb5;
frames[14][26][34] = 8'hb1;
frames[14][26][35] = 8'hb5;
frames[14][26][36] = 8'hd6;
frames[14][26][37] = 8'hb6;
frames[14][26][38] = 8'hb5;
frames[14][26][39] = 8'hb5;
frames[14][27][0] = 8'h44;
frames[14][27][1] = 8'h44;
frames[14][27][2] = 8'h24;
frames[14][27][3] = 8'h24;
frames[14][27][4] = 8'h24;
frames[14][27][5] = 8'h24;
frames[14][27][6] = 8'h24;
frames[14][27][7] = 8'h44;
frames[14][27][8] = 8'h24;
frames[14][27][9] = 8'h24;
frames[14][27][10] = 8'h20;
frames[14][27][11] = 8'h24;
frames[14][27][12] = 8'h44;
frames[14][27][13] = 8'h44;
frames[14][27][14] = 8'h64;
frames[14][27][15] = 8'h64;
frames[14][27][16] = 8'h68;
frames[14][27][17] = 8'h68;
frames[14][27][18] = 8'h68;
frames[14][27][19] = 8'h8d;
frames[14][27][20] = 8'hb1;
frames[14][27][21] = 8'hd1;
frames[14][27][22] = 8'hd1;
frames[14][27][23] = 8'hd6;
frames[14][27][24] = 8'hd5;
frames[14][27][25] = 8'hb1;
frames[14][27][26] = 8'hb1;
frames[14][27][27] = 8'hb5;
frames[14][27][28] = 8'hb5;
frames[14][27][29] = 8'hb1;
frames[14][27][30] = 8'hb1;
frames[14][27][31] = 8'hb5;
frames[14][27][32] = 8'hb5;
frames[14][27][33] = 8'hb1;
frames[14][27][34] = 8'hb1;
frames[14][27][35] = 8'hb5;
frames[14][27][36] = 8'hb5;
frames[14][27][37] = 8'hb1;
frames[14][27][38] = 8'hb1;
frames[14][27][39] = 8'hb1;
frames[14][28][0] = 8'h44;
frames[14][28][1] = 8'h44;
frames[14][28][2] = 8'h44;
frames[14][28][3] = 8'h44;
frames[14][28][4] = 8'h44;
frames[14][28][5] = 8'h44;
frames[14][28][6] = 8'h44;
frames[14][28][7] = 8'h44;
frames[14][28][8] = 8'h44;
frames[14][28][9] = 8'h44;
frames[14][28][10] = 8'h44;
frames[14][28][11] = 8'h44;
frames[14][28][12] = 8'h44;
frames[14][28][13] = 8'h68;
frames[14][28][14] = 8'h68;
frames[14][28][15] = 8'h68;
frames[14][28][16] = 8'h8c;
frames[14][28][17] = 8'hb1;
frames[14][28][18] = 8'hd2;
frames[14][28][19] = 8'hd6;
frames[14][28][20] = 8'hd6;
frames[14][28][21] = 8'hd6;
frames[14][28][22] = 8'hd6;
frames[14][28][23] = 8'hd6;
frames[14][28][24] = 8'hd1;
frames[14][28][25] = 8'hd6;
frames[14][28][26] = 8'hb1;
frames[14][28][27] = 8'hb1;
frames[14][28][28] = 8'hd6;
frames[14][28][29] = 8'hb1;
frames[14][28][30] = 8'hb1;
frames[14][28][31] = 8'hb5;
frames[14][28][32] = 8'hd5;
frames[14][28][33] = 8'hb5;
frames[14][28][34] = 8'hb5;
frames[14][28][35] = 8'hb1;
frames[14][28][36] = 8'hb1;
frames[14][28][37] = 8'hb1;
frames[14][28][38] = 8'h91;
frames[14][28][39] = 8'h91;
frames[14][29][0] = 8'h68;
frames[14][29][1] = 8'h64;
frames[14][29][2] = 8'h44;
frames[14][29][3] = 8'h44;
frames[14][29][4] = 8'h44;
frames[14][29][5] = 8'h44;
frames[14][29][6] = 8'h44;
frames[14][29][7] = 8'h44;
frames[14][29][8] = 8'h44;
frames[14][29][9] = 8'h44;
frames[14][29][10] = 8'h44;
frames[14][29][11] = 8'h44;
frames[14][29][12] = 8'h68;
frames[14][29][13] = 8'h68;
frames[14][29][14] = 8'h88;
frames[14][29][15] = 8'hb1;
frames[14][29][16] = 8'hd6;
frames[14][29][17] = 8'hfa;
frames[14][29][18] = 8'hd6;
frames[14][29][19] = 8'hd6;
frames[14][29][20] = 8'hd6;
frames[14][29][21] = 8'hd6;
frames[14][29][22] = 8'hd6;
frames[14][29][23] = 8'hd6;
frames[14][29][24] = 8'hb1;
frames[14][29][25] = 8'hb1;
frames[14][29][26] = 8'hb1;
frames[14][29][27] = 8'had;
frames[14][29][28] = 8'hd5;
frames[14][29][29] = 8'hb1;
frames[14][29][30] = 8'hb1;
frames[14][29][31] = 8'hb1;
frames[14][29][32] = 8'hb1;
frames[14][29][33] = 8'hb1;
frames[14][29][34] = 8'hb5;
frames[14][29][35] = 8'hb1;
frames[14][29][36] = 8'h91;
frames[14][29][37] = 8'h91;
frames[14][29][38] = 8'h8d;
frames[14][29][39] = 8'h8d;
frames[15][0][0] = 8'h89;
frames[15][0][1] = 8'h89;
frames[15][0][2] = 8'h89;
frames[15][0][3] = 8'h89;
frames[15][0][4] = 8'h89;
frames[15][0][5] = 8'h89;
frames[15][0][6] = 8'h00;
frames[15][0][7] = 8'h00;
frames[15][0][8] = 8'h00;
frames[15][0][9] = 8'h00;
frames[15][0][10] = 8'h00;
frames[15][0][11] = 8'h00;
frames[15][0][12] = 8'h00;
frames[15][0][13] = 8'h00;
frames[15][0][14] = 8'h00;
frames[15][0][15] = 8'h00;
frames[15][0][16] = 8'h00;
frames[15][0][17] = 8'h00;
frames[15][0][18] = 8'h00;
frames[15][0][19] = 8'h00;
frames[15][0][20] = 8'h00;
frames[15][0][21] = 8'h00;
frames[15][0][22] = 8'h00;
frames[15][0][23] = 8'h00;
frames[15][0][24] = 8'h20;
frames[15][0][25] = 8'h8d;
frames[15][0][26] = 8'h89;
frames[15][0][27] = 8'h64;
frames[15][0][28] = 8'h89;
frames[15][0][29] = 8'had;
frames[15][0][30] = 8'ha9;
frames[15][0][31] = 8'ha9;
frames[15][0][32] = 8'h8d;
frames[15][0][33] = 8'h44;
frames[15][0][34] = 8'h8d;
frames[15][0][35] = 8'hda;
frames[15][0][36] = 8'hd6;
frames[15][0][37] = 8'hfb;
frames[15][0][38] = 8'hdb;
frames[15][0][39] = 8'hda;
frames[15][1][0] = 8'h88;
frames[15][1][1] = 8'h88;
frames[15][1][2] = 8'h88;
frames[15][1][3] = 8'h88;
frames[15][1][4] = 8'h88;
frames[15][1][5] = 8'h89;
frames[15][1][6] = 8'h24;
frames[15][1][7] = 8'h00;
frames[15][1][8] = 8'h00;
frames[15][1][9] = 8'h00;
frames[15][1][10] = 8'h00;
frames[15][1][11] = 8'h00;
frames[15][1][12] = 8'h00;
frames[15][1][13] = 8'h00;
frames[15][1][14] = 8'h00;
frames[15][1][15] = 8'h00;
frames[15][1][16] = 8'h00;
frames[15][1][17] = 8'h00;
frames[15][1][18] = 8'h00;
frames[15][1][19] = 8'h00;
frames[15][1][20] = 8'h00;
frames[15][1][21] = 8'h00;
frames[15][1][22] = 8'h00;
frames[15][1][23] = 8'h00;
frames[15][1][24] = 8'h40;
frames[15][1][25] = 8'h8d;
frames[15][1][26] = 8'h88;
frames[15][1][27] = 8'h64;
frames[15][1][28] = 8'had;
frames[15][1][29] = 8'had;
frames[15][1][30] = 8'ha9;
frames[15][1][31] = 8'ha9;
frames[15][1][32] = 8'h8d;
frames[15][1][33] = 8'h40;
frames[15][1][34] = 8'h69;
frames[15][1][35] = 8'hda;
frames[15][1][36] = 8'hdb;
frames[15][1][37] = 8'hfb;
frames[15][1][38] = 8'hdb;
frames[15][1][39] = 8'hdb;
frames[15][2][0] = 8'h88;
frames[15][2][1] = 8'h89;
frames[15][2][2] = 8'h64;
frames[15][2][3] = 8'h64;
frames[15][2][4] = 8'h64;
frames[15][2][5] = 8'h89;
frames[15][2][6] = 8'h44;
frames[15][2][7] = 8'h00;
frames[15][2][8] = 8'h00;
frames[15][2][9] = 8'h00;
frames[15][2][10] = 8'h00;
frames[15][2][11] = 8'h00;
frames[15][2][12] = 8'h00;
frames[15][2][13] = 8'h00;
frames[15][2][14] = 8'h00;
frames[15][2][15] = 8'h00;
frames[15][2][16] = 8'h00;
frames[15][2][17] = 8'h00;
frames[15][2][18] = 8'h00;
frames[15][2][19] = 8'h00;
frames[15][2][20] = 8'h00;
frames[15][2][21] = 8'h00;
frames[15][2][22] = 8'h00;
frames[15][2][23] = 8'h00;
frames[15][2][24] = 8'h44;
frames[15][2][25] = 8'h8d;
frames[15][2][26] = 8'h64;
frames[15][2][27] = 8'h88;
frames[15][2][28] = 8'had;
frames[15][2][29] = 8'had;
frames[15][2][30] = 8'h89;
frames[15][2][31] = 8'had;
frames[15][2][32] = 8'h8d;
frames[15][2][33] = 8'h20;
frames[15][2][34] = 8'h48;
frames[15][2][35] = 8'hda;
frames[15][2][36] = 8'hfb;
frames[15][2][37] = 8'hdb;
frames[15][2][38] = 8'h4d;
frames[15][2][39] = 8'hbb;
frames[15][3][0] = 8'h88;
frames[15][3][1] = 8'h89;
frames[15][3][2] = 8'h68;
frames[15][3][3] = 8'h20;
frames[15][3][4] = 8'h40;
frames[15][3][5] = 8'h68;
frames[15][3][6] = 8'h69;
frames[15][3][7] = 8'h20;
frames[15][3][8] = 8'h00;
frames[15][3][9] = 8'h00;
frames[15][3][10] = 8'h00;
frames[15][3][11] = 8'h00;
frames[15][3][12] = 8'h00;
frames[15][3][13] = 8'h00;
frames[15][3][14] = 8'h00;
frames[15][3][15] = 8'h20;
frames[15][3][16] = 8'h24;
frames[15][3][17] = 8'h24;
frames[15][3][18] = 8'h24;
frames[15][3][19] = 8'h48;
frames[15][3][20] = 8'h48;
frames[15][3][21] = 8'h44;
frames[15][3][22] = 8'h24;
frames[15][3][23] = 8'h00;
frames[15][3][24] = 8'h68;
frames[15][3][25] = 8'h89;
frames[15][3][26] = 8'h64;
frames[15][3][27] = 8'had;
frames[15][3][28] = 8'had;
frames[15][3][29] = 8'h89;
frames[15][3][30] = 8'h8d;
frames[15][3][31] = 8'had;
frames[15][3][32] = 8'h44;
frames[15][3][33] = 8'h00;
frames[15][3][34] = 8'h24;
frames[15][3][35] = 8'hda;
frames[15][3][36] = 8'hdb;
frames[15][3][37] = 8'hda;
frames[15][3][38] = 8'h49;
frames[15][3][39] = 8'hb7;
frames[15][4][0] = 8'h68;
frames[15][4][1] = 8'h89;
frames[15][4][2] = 8'h89;
frames[15][4][3] = 8'h40;
frames[15][4][4] = 8'h20;
frames[15][4][5] = 8'h44;
frames[15][4][6] = 8'h89;
frames[15][4][7] = 8'h44;
frames[15][4][8] = 8'h00;
frames[15][4][9] = 8'h24;
frames[15][4][10] = 8'h44;
frames[15][4][11] = 8'h69;
frames[15][4][12] = 8'h6d;
frames[15][4][13] = 8'h8d;
frames[15][4][14] = 8'h8d;
frames[15][4][15] = 8'h8d;
frames[15][4][16] = 8'h91;
frames[15][4][17] = 8'hb1;
frames[15][4][18] = 8'hb1;
frames[15][4][19] = 8'hb5;
frames[15][4][20] = 8'hd6;
frames[15][4][21] = 8'hd6;
frames[15][4][22] = 8'hb2;
frames[15][4][23] = 8'h8d;
frames[15][4][24] = 8'h89;
frames[15][4][25] = 8'h64;
frames[15][4][26] = 8'h89;
frames[15][4][27] = 8'had;
frames[15][4][28] = 8'h89;
frames[15][4][29] = 8'h88;
frames[15][4][30] = 8'had;
frames[15][4][31] = 8'h89;
frames[15][4][32] = 8'h00;
frames[15][4][33] = 8'h00;
frames[15][4][34] = 8'h20;
frames[15][4][35] = 8'hb6;
frames[15][4][36] = 8'hfb;
frames[15][4][37] = 8'hda;
frames[15][4][38] = 8'h92;
frames[15][4][39] = 8'hdb;
frames[15][5][0] = 8'h88;
frames[15][5][1] = 8'h64;
frames[15][5][2] = 8'h89;
frames[15][5][3] = 8'h68;
frames[15][5][4] = 8'h20;
frames[15][5][5] = 8'h20;
frames[15][5][6] = 8'h68;
frames[15][5][7] = 8'h88;
frames[15][5][8] = 8'h8d;
frames[15][5][9] = 8'h8d;
frames[15][5][10] = 8'hb1;
frames[15][5][11] = 8'hb1;
frames[15][5][12] = 8'hb1;
frames[15][5][13] = 8'hb1;
frames[15][5][14] = 8'hb1;
frames[15][5][15] = 8'hb1;
frames[15][5][16] = 8'hb1;
frames[15][5][17] = 8'hb1;
frames[15][5][18] = 8'hb1;
frames[15][5][19] = 8'hb1;
frames[15][5][20] = 8'hb1;
frames[15][5][21] = 8'hd5;
frames[15][5][22] = 8'hd6;
frames[15][5][23] = 8'hb1;
frames[15][5][24] = 8'h89;
frames[15][5][25] = 8'h89;
frames[15][5][26] = 8'had;
frames[15][5][27] = 8'h89;
frames[15][5][28] = 8'h88;
frames[15][5][29] = 8'had;
frames[15][5][30] = 8'h8d;
frames[15][5][31] = 8'h44;
frames[15][5][32] = 8'h00;
frames[15][5][33] = 8'h00;
frames[15][5][34] = 8'h00;
frames[15][5][35] = 8'hb6;
frames[15][5][36] = 8'hfb;
frames[15][5][37] = 8'hff;
frames[15][5][38] = 8'hff;
frames[15][5][39] = 8'hdb;
frames[15][6][0] = 8'h88;
frames[15][6][1] = 8'h64;
frames[15][6][2] = 8'h84;
frames[15][6][3] = 8'h89;
frames[15][6][4] = 8'h89;
frames[15][6][5] = 8'h64;
frames[15][6][6] = 8'h88;
frames[15][6][7] = 8'h88;
frames[15][6][8] = 8'h89;
frames[15][6][9] = 8'h8d;
frames[15][6][10] = 8'h8d;
frames[15][6][11] = 8'h8d;
frames[15][6][12] = 8'h8d;
frames[15][6][13] = 8'h8d;
frames[15][6][14] = 8'h8d;
frames[15][6][15] = 8'hb1;
frames[15][6][16] = 8'hb1;
frames[15][6][17] = 8'hb1;
frames[15][6][18] = 8'hb1;
frames[15][6][19] = 8'hb1;
frames[15][6][20] = 8'hb1;
frames[15][6][21] = 8'hb1;
frames[15][6][22] = 8'hb1;
frames[15][6][23] = 8'had;
frames[15][6][24] = 8'h89;
frames[15][6][25] = 8'had;
frames[15][6][26] = 8'h89;
frames[15][6][27] = 8'h68;
frames[15][6][28] = 8'h89;
frames[15][6][29] = 8'had;
frames[15][6][30] = 8'h69;
frames[15][6][31] = 8'h20;
frames[15][6][32] = 8'h00;
frames[15][6][33] = 8'h00;
frames[15][6][34] = 8'h00;
frames[15][6][35] = 8'hb6;
frames[15][6][36] = 8'hdb;
frames[15][6][37] = 8'hda;
frames[15][6][38] = 8'hda;
frames[15][6][39] = 8'hda;
frames[15][7][0] = 8'h64;
frames[15][7][1] = 8'h89;
frames[15][7][2] = 8'h88;
frames[15][7][3] = 8'h88;
frames[15][7][4] = 8'h88;
frames[15][7][5] = 8'h64;
frames[15][7][6] = 8'h8d;
frames[15][7][7] = 8'h8d;
frames[15][7][8] = 8'h89;
frames[15][7][9] = 8'h8d;
frames[15][7][10] = 8'h8d;
frames[15][7][11] = 8'h8d;
frames[15][7][12] = 8'h8d;
frames[15][7][13] = 8'h8d;
frames[15][7][14] = 8'h8d;
frames[15][7][15] = 8'hb1;
frames[15][7][16] = 8'hb1;
frames[15][7][17] = 8'hb1;
frames[15][7][18] = 8'hb1;
frames[15][7][19] = 8'hb1;
frames[15][7][20] = 8'hb1;
frames[15][7][21] = 8'hb1;
frames[15][7][22] = 8'hb1;
frames[15][7][23] = 8'had;
frames[15][7][24] = 8'ha9;
frames[15][7][25] = 8'h89;
frames[15][7][26] = 8'h89;
frames[15][7][27] = 8'h89;
frames[15][7][28] = 8'had;
frames[15][7][29] = 8'h89;
frames[15][7][30] = 8'h44;
frames[15][7][31] = 8'h20;
frames[15][7][32] = 8'h00;
frames[15][7][33] = 8'h00;
frames[15][7][34] = 8'h48;
frames[15][7][35] = 8'hb6;
frames[15][7][36] = 8'hfb;
frames[15][7][37] = 8'hdb;
frames[15][7][38] = 8'hda;
frames[15][7][39] = 8'hb6;
frames[15][8][0] = 8'h20;
frames[15][8][1] = 8'h68;
frames[15][8][2] = 8'h89;
frames[15][8][3] = 8'h89;
frames[15][8][4] = 8'h88;
frames[15][8][5] = 8'h64;
frames[15][8][6] = 8'h44;
frames[15][8][7] = 8'had;
frames[15][8][8] = 8'hb1;
frames[15][8][9] = 8'h8d;
frames[15][8][10] = 8'h8d;
frames[15][8][11] = 8'h8d;
frames[15][8][12] = 8'h8d;
frames[15][8][13] = 8'h8d;
frames[15][8][14] = 8'h8d;
frames[15][8][15] = 8'hb1;
frames[15][8][16] = 8'hb1;
frames[15][8][17] = 8'hb1;
frames[15][8][18] = 8'hb1;
frames[15][8][19] = 8'hb1;
frames[15][8][20] = 8'hb1;
frames[15][8][21] = 8'hb1;
frames[15][8][22] = 8'h8d;
frames[15][8][23] = 8'h68;
frames[15][8][24] = 8'h68;
frames[15][8][25] = 8'h64;
frames[15][8][26] = 8'h89;
frames[15][8][27] = 8'h89;
frames[15][8][28] = 8'h48;
frames[15][8][29] = 8'h44;
frames[15][8][30] = 8'h24;
frames[15][8][31] = 8'h24;
frames[15][8][32] = 8'h24;
frames[15][8][33] = 8'h49;
frames[15][8][34] = 8'hdb;
frames[15][8][35] = 8'hff;
frames[15][8][36] = 8'hff;
frames[15][8][37] = 8'hfb;
frames[15][8][38] = 8'hda;
frames[15][8][39] = 8'hb2;
frames[15][9][0] = 8'h24;
frames[15][9][1] = 8'h24;
frames[15][9][2] = 8'h44;
frames[15][9][3] = 8'h44;
frames[15][9][4] = 8'h64;
frames[15][9][5] = 8'h44;
frames[15][9][6] = 8'h20;
frames[15][9][7] = 8'h44;
frames[15][9][8] = 8'h8d;
frames[15][9][9] = 8'hb1;
frames[15][9][10] = 8'hb1;
frames[15][9][11] = 8'hb1;
frames[15][9][12] = 8'hb1;
frames[15][9][13] = 8'hb1;
frames[15][9][14] = 8'hb1;
frames[15][9][15] = 8'hb1;
frames[15][9][16] = 8'hb1;
frames[15][9][17] = 8'hb1;
frames[15][9][18] = 8'hb1;
frames[15][9][19] = 8'hb1;
frames[15][9][20] = 8'hb1;
frames[15][9][21] = 8'hb1;
frames[15][9][22] = 8'h69;
frames[15][9][23] = 8'h44;
frames[15][9][24] = 8'h44;
frames[15][9][25] = 8'h44;
frames[15][9][26] = 8'h44;
frames[15][9][27] = 8'h24;
frames[15][9][28] = 8'h24;
frames[15][9][29] = 8'h20;
frames[15][9][30] = 8'h24;
frames[15][9][31] = 8'h24;
frames[15][9][32] = 8'h44;
frames[15][9][33] = 8'h8d;
frames[15][9][34] = 8'hdb;
frames[15][9][35] = 8'hfb;
frames[15][9][36] = 8'hff;
frames[15][9][37] = 8'hdb;
frames[15][9][38] = 8'hda;
frames[15][9][39] = 8'h91;
frames[15][10][0] = 8'h49;
frames[15][10][1] = 8'h24;
frames[15][10][2] = 8'h00;
frames[15][10][3] = 8'h20;
frames[15][10][4] = 8'h20;
frames[15][10][5] = 8'h20;
frames[15][10][6] = 8'h20;
frames[15][10][7] = 8'h20;
frames[15][10][8] = 8'h44;
frames[15][10][9] = 8'h8d;
frames[15][10][10] = 8'hb1;
frames[15][10][11] = 8'hb2;
frames[15][10][12] = 8'hb1;
frames[15][10][13] = 8'hb1;
frames[15][10][14] = 8'hb1;
frames[15][10][15] = 8'hb1;
frames[15][10][16] = 8'hd6;
frames[15][10][17] = 8'hd6;
frames[15][10][18] = 8'hd5;
frames[15][10][19] = 8'hd5;
frames[15][10][20] = 8'hb1;
frames[15][10][21] = 8'hb1;
frames[15][10][22] = 8'hb1;
frames[15][10][23] = 8'h8d;
frames[15][10][24] = 8'h6d;
frames[15][10][25] = 8'h68;
frames[15][10][26] = 8'h24;
frames[15][10][27] = 8'h24;
frames[15][10][28] = 8'h24;
frames[15][10][29] = 8'h24;
frames[15][10][30] = 8'h24;
frames[15][10][31] = 8'h24;
frames[15][10][32] = 8'h48;
frames[15][10][33] = 8'h92;
frames[15][10][34] = 8'hdb;
frames[15][10][35] = 8'hfb;
frames[15][10][36] = 8'hdb;
frames[15][10][37] = 8'hdb;
frames[15][10][38] = 8'hda;
frames[15][10][39] = 8'h91;
frames[15][11][0] = 8'h49;
frames[15][11][1] = 8'h24;
frames[15][11][2] = 8'h20;
frames[15][11][3] = 8'h00;
frames[15][11][4] = 8'h24;
frames[15][11][5] = 8'h48;
frames[15][11][6] = 8'h68;
frames[15][11][7] = 8'h69;
frames[15][11][8] = 8'h8d;
frames[15][11][9] = 8'h68;
frames[15][11][10] = 8'h68;
frames[15][11][11] = 8'h8d;
frames[15][11][12] = 8'h8d;
frames[15][11][13] = 8'hb1;
frames[15][11][14] = 8'hb1;
frames[15][11][15] = 8'hb1;
frames[15][11][16] = 8'hd5;
frames[15][11][17] = 8'hd5;
frames[15][11][18] = 8'hd6;
frames[15][11][19] = 8'hd6;
frames[15][11][20] = 8'hb6;
frames[15][11][21] = 8'hb1;
frames[15][11][22] = 8'hb1;
frames[15][11][23] = 8'hb1;
frames[15][11][24] = 8'hb1;
frames[15][11][25] = 8'h8d;
frames[15][11][26] = 8'h44;
frames[15][11][27] = 8'h20;
frames[15][11][28] = 8'h20;
frames[15][11][29] = 8'h20;
frames[15][11][30] = 8'h20;
frames[15][11][31] = 8'h20;
frames[15][11][32] = 8'h48;
frames[15][11][33] = 8'hb2;
frames[15][11][34] = 8'hdb;
frames[15][11][35] = 8'hdb;
frames[15][11][36] = 8'hdb;
frames[15][11][37] = 8'hdb;
frames[15][11][38] = 8'hda;
frames[15][11][39] = 8'h91;
frames[15][12][0] = 8'h49;
frames[15][12][1] = 8'h24;
frames[15][12][2] = 8'h24;
frames[15][12][3] = 8'h24;
frames[15][12][4] = 8'h8d;
frames[15][12][5] = 8'h8d;
frames[15][12][6] = 8'h8d;
frames[15][12][7] = 8'hb1;
frames[15][12][8] = 8'had;
frames[15][12][9] = 8'h8c;
frames[15][12][10] = 8'h68;
frames[15][12][11] = 8'h8d;
frames[15][12][12] = 8'h68;
frames[15][12][13] = 8'h8d;
frames[15][12][14] = 8'hb1;
frames[15][12][15] = 8'hb1;
frames[15][12][16] = 8'hb5;
frames[15][12][17] = 8'hd5;
frames[15][12][18] = 8'hd6;
frames[15][12][19] = 8'hb5;
frames[15][12][20] = 8'h91;
frames[15][12][21] = 8'hb1;
frames[15][12][22] = 8'hb1;
frames[15][12][23] = 8'hb1;
frames[15][12][24] = 8'h8d;
frames[15][12][25] = 8'h48;
frames[15][12][26] = 8'h20;
frames[15][12][27] = 8'h20;
frames[15][12][28] = 8'h20;
frames[15][12][29] = 8'h20;
frames[15][12][30] = 8'h20;
frames[15][12][31] = 8'h00;
frames[15][12][32] = 8'h44;
frames[15][12][33] = 8'hb6;
frames[15][12][34] = 8'hdb;
frames[15][12][35] = 8'hdb;
frames[15][12][36] = 8'hdb;
frames[15][12][37] = 8'hdb;
frames[15][12][38] = 8'hd6;
frames[15][12][39] = 8'hb6;
frames[15][13][0] = 8'h48;
frames[15][13][1] = 8'h24;
frames[15][13][2] = 8'h24;
frames[15][13][3] = 8'h6d;
frames[15][13][4] = 8'h91;
frames[15][13][5] = 8'h91;
frames[15][13][6] = 8'h8d;
frames[15][13][7] = 8'hd5;
frames[15][13][8] = 8'hb1;
frames[15][13][9] = 8'hb1;
frames[15][13][10] = 8'h8c;
frames[15][13][11] = 8'hb1;
frames[15][13][12] = 8'hb1;
frames[15][13][13] = 8'hb1;
frames[15][13][14] = 8'hb1;
frames[15][13][15] = 8'hb1;
frames[15][13][16] = 8'hb1;
frames[15][13][17] = 8'hb1;
frames[15][13][18] = 8'hb1;
frames[15][13][19] = 8'hb1;
frames[15][13][20] = 8'hb1;
frames[15][13][21] = 8'hd5;
frames[15][13][22] = 8'hb1;
frames[15][13][23] = 8'h8d;
frames[15][13][24] = 8'h48;
frames[15][13][25] = 8'h24;
frames[15][13][26] = 8'h20;
frames[15][13][27] = 8'h20;
frames[15][13][28] = 8'h20;
frames[15][13][29] = 8'h20;
frames[15][13][30] = 8'h00;
frames[15][13][31] = 8'h00;
frames[15][13][32] = 8'h24;
frames[15][13][33] = 8'h92;
frames[15][13][34] = 8'hdb;
frames[15][13][35] = 8'hdb;
frames[15][13][36] = 8'hdb;
frames[15][13][37] = 8'hdb;
frames[15][13][38] = 8'hd6;
frames[15][13][39] = 8'hb6;
frames[15][14][0] = 8'h24;
frames[15][14][1] = 8'h24;
frames[15][14][2] = 8'h24;
frames[15][14][3] = 8'h24;
frames[15][14][4] = 8'h6d;
frames[15][14][5] = 8'hb6;
frames[15][14][6] = 8'hd5;
frames[15][14][7] = 8'hd5;
frames[15][14][8] = 8'hb1;
frames[15][14][9] = 8'hd5;
frames[15][14][10] = 8'hb1;
frames[15][14][11] = 8'hd6;
frames[15][14][12] = 8'hd6;
frames[15][14][13] = 8'hd6;
frames[15][14][14] = 8'hd6;
frames[15][14][15] = 8'hb5;
frames[15][14][16] = 8'hd5;
frames[15][14][17] = 8'had;
frames[15][14][18] = 8'h68;
frames[15][14][19] = 8'had;
frames[15][14][20] = 8'hb2;
frames[15][14][21] = 8'hb1;
frames[15][14][22] = 8'h69;
frames[15][14][23] = 8'h44;
frames[15][14][24] = 8'h24;
frames[15][14][25] = 8'h24;
frames[15][14][26] = 8'h24;
frames[15][14][27] = 8'h20;
frames[15][14][28] = 8'h20;
frames[15][14][29] = 8'h20;
frames[15][14][30] = 8'h20;
frames[15][14][31] = 8'h00;
frames[15][14][32] = 8'h24;
frames[15][14][33] = 8'h92;
frames[15][14][34] = 8'hfb;
frames[15][14][35] = 8'hdb;
frames[15][14][36] = 8'hdb;
frames[15][14][37] = 8'hdb;
frames[15][14][38] = 8'hd6;
frames[15][14][39] = 8'hb6;
frames[15][15][0] = 8'h24;
frames[15][15][1] = 8'h24;
frames[15][15][2] = 8'h48;
frames[15][15][3] = 8'h24;
frames[15][15][4] = 8'h44;
frames[15][15][5] = 8'h48;
frames[15][15][6] = 8'hb1;
frames[15][15][7] = 8'hd6;
frames[15][15][8] = 8'hd5;
frames[15][15][9] = 8'hd5;
frames[15][15][10] = 8'hd6;
frames[15][15][11] = 8'hd6;
frames[15][15][12] = 8'hd6;
frames[15][15][13] = 8'hd6;
frames[15][15][14] = 8'hd6;
frames[15][15][15] = 8'hd5;
frames[15][15][16] = 8'hb5;
frames[15][15][17] = 8'hb5;
frames[15][15][18] = 8'hb1;
frames[15][15][19] = 8'h8d;
frames[15][15][20] = 8'h44;
frames[15][15][21] = 8'h24;
frames[15][15][22] = 8'h24;
frames[15][15][23] = 8'h24;
frames[15][15][24] = 8'h24;
frames[15][15][25] = 8'h24;
frames[15][15][26] = 8'h24;
frames[15][15][27] = 8'h20;
frames[15][15][28] = 8'h20;
frames[15][15][29] = 8'h20;
frames[15][15][30] = 8'h24;
frames[15][15][31] = 8'h20;
frames[15][15][32] = 8'h24;
frames[15][15][33] = 8'h6d;
frames[15][15][34] = 8'hfb;
frames[15][15][35] = 8'hdb;
frames[15][15][36] = 8'hdb;
frames[15][15][37] = 8'hdb;
frames[15][15][38] = 8'hd6;
frames[15][15][39] = 8'hb6;
frames[15][16][0] = 8'h24;
frames[15][16][1] = 8'h24;
frames[15][16][2] = 8'h48;
frames[15][16][3] = 8'h44;
frames[15][16][4] = 8'h44;
frames[15][16][5] = 8'h44;
frames[15][16][6] = 8'h44;
frames[15][16][7] = 8'h48;
frames[15][16][8] = 8'h8d;
frames[15][16][9] = 8'h68;
frames[15][16][10] = 8'hb6;
frames[15][16][11] = 8'hd6;
frames[15][16][12] = 8'hd6;
frames[15][16][13] = 8'hb6;
frames[15][16][14] = 8'hd6;
frames[15][16][15] = 8'hd6;
frames[15][16][16] = 8'hd6;
frames[15][16][17] = 8'hd6;
frames[15][16][18] = 8'hd6;
frames[15][16][19] = 8'hb1;
frames[15][16][20] = 8'h6d;
frames[15][16][21] = 8'h44;
frames[15][16][22] = 8'h24;
frames[15][16][23] = 8'h24;
frames[15][16][24] = 8'h24;
frames[15][16][25] = 8'h24;
frames[15][16][26] = 8'h24;
frames[15][16][27] = 8'h24;
frames[15][16][28] = 8'h24;
frames[15][16][29] = 8'h24;
frames[15][16][30] = 8'h24;
frames[15][16][31] = 8'h24;
frames[15][16][32] = 8'h24;
frames[15][16][33] = 8'h49;
frames[15][16][34] = 8'hdb;
frames[15][16][35] = 8'hfb;
frames[15][16][36] = 8'hdb;
frames[15][16][37] = 8'hdb;
frames[15][16][38] = 8'hd6;
frames[15][16][39] = 8'hb6;
frames[15][17][0] = 8'h24;
frames[15][17][1] = 8'h24;
frames[15][17][2] = 8'h49;
frames[15][17][3] = 8'h44;
frames[15][17][4] = 8'h24;
frames[15][17][5] = 8'h24;
frames[15][17][6] = 8'h44;
frames[15][17][7] = 8'h69;
frames[15][17][8] = 8'hb6;
frames[15][17][9] = 8'hb1;
frames[15][17][10] = 8'hd6;
frames[15][17][11] = 8'hda;
frames[15][17][12] = 8'hda;
frames[15][17][13] = 8'hd6;
frames[15][17][14] = 8'hd6;
frames[15][17][15] = 8'hd6;
frames[15][17][16] = 8'hd6;
frames[15][17][17] = 8'hda;
frames[15][17][18] = 8'hd6;
frames[15][17][19] = 8'hda;
frames[15][17][20] = 8'hd6;
frames[15][17][21] = 8'hb1;
frames[15][17][22] = 8'h8d;
frames[15][17][23] = 8'h44;
frames[15][17][24] = 8'h24;
frames[15][17][25] = 8'h24;
frames[15][17][26] = 8'h24;
frames[15][17][27] = 8'h24;
frames[15][17][28] = 8'h24;
frames[15][17][29] = 8'h24;
frames[15][17][30] = 8'h44;
frames[15][17][31] = 8'h44;
frames[15][17][32] = 8'h24;
frames[15][17][33] = 8'h44;
frames[15][17][34] = 8'hb6;
frames[15][17][35] = 8'hfb;
frames[15][17][36] = 8'hdb;
frames[15][17][37] = 8'hda;
frames[15][17][38] = 8'hd6;
frames[15][17][39] = 8'hb6;
frames[15][18][0] = 8'h24;
frames[15][18][1] = 8'h44;
frames[15][18][2] = 8'h48;
frames[15][18][3] = 8'h24;
frames[15][18][4] = 8'h44;
frames[15][18][5] = 8'h6d;
frames[15][18][6] = 8'had;
frames[15][18][7] = 8'hb1;
frames[15][18][8] = 8'had;
frames[15][18][9] = 8'had;
frames[15][18][10] = 8'hd6;
frames[15][18][11] = 8'hd6;
frames[15][18][12] = 8'hd6;
frames[15][18][13] = 8'hd6;
frames[15][18][14] = 8'hd6;
frames[15][18][15] = 8'hd6;
frames[15][18][16] = 8'hda;
frames[15][18][17] = 8'hda;
frames[15][18][18] = 8'hd6;
frames[15][18][19] = 8'hd6;
frames[15][18][20] = 8'hd6;
frames[15][18][21] = 8'hb6;
frames[15][18][22] = 8'hb1;
frames[15][18][23] = 8'hb1;
frames[15][18][24] = 8'h6d;
frames[15][18][25] = 8'h24;
frames[15][18][26] = 8'h24;
frames[15][18][27] = 8'h24;
frames[15][18][28] = 8'h24;
frames[15][18][29] = 8'h24;
frames[15][18][30] = 8'h44;
frames[15][18][31] = 8'h48;
frames[15][18][32] = 8'h44;
frames[15][18][33] = 8'h44;
frames[15][18][34] = 8'h91;
frames[15][18][35] = 8'hfb;
frames[15][18][36] = 8'hdb;
frames[15][18][37] = 8'hda;
frames[15][18][38] = 8'hd6;
frames[15][18][39] = 8'hd6;
frames[15][19][0] = 8'h24;
frames[15][19][1] = 8'h49;
frames[15][19][2] = 8'h48;
frames[15][19][3] = 8'h48;
frames[15][19][4] = 8'h8d;
frames[15][19][5] = 8'hd6;
frames[15][19][6] = 8'hb1;
frames[15][19][7] = 8'h8d;
frames[15][19][8] = 8'had;
frames[15][19][9] = 8'hd1;
frames[15][19][10] = 8'hd6;
frames[15][19][11] = 8'hd6;
frames[15][19][12] = 8'hd5;
frames[15][19][13] = 8'hd5;
frames[15][19][14] = 8'hd6;
frames[15][19][15] = 8'hd6;
frames[15][19][16] = 8'hd6;
frames[15][19][17] = 8'hd6;
frames[15][19][18] = 8'hd5;
frames[15][19][19] = 8'hb1;
frames[15][19][20] = 8'hd5;
frames[15][19][21] = 8'hb5;
frames[15][19][22] = 8'hd6;
frames[15][19][23] = 8'hb5;
frames[15][19][24] = 8'hb6;
frames[15][19][25] = 8'h91;
frames[15][19][26] = 8'h69;
frames[15][19][27] = 8'h44;
frames[15][19][28] = 8'h24;
frames[15][19][29] = 8'h44;
frames[15][19][30] = 8'h48;
frames[15][19][31] = 8'h49;
frames[15][19][32] = 8'h44;
frames[15][19][33] = 8'h44;
frames[15][19][34] = 8'h6d;
frames[15][19][35] = 8'hdb;
frames[15][19][36] = 8'hdb;
frames[15][19][37] = 8'hda;
frames[15][19][38] = 8'hd6;
frames[15][19][39] = 8'hd6;
frames[15][20][0] = 8'h24;
frames[15][20][1] = 8'h49;
frames[15][20][2] = 8'h44;
frames[15][20][3] = 8'h6d;
frames[15][20][4] = 8'hb6;
frames[15][20][5] = 8'hd6;
frames[15][20][6] = 8'hb1;
frames[15][20][7] = 8'hb1;
frames[15][20][8] = 8'h8d;
frames[15][20][9] = 8'hd1;
frames[15][20][10] = 8'hd6;
frames[15][20][11] = 8'hd6;
frames[15][20][12] = 8'hd5;
frames[15][20][13] = 8'hb5;
frames[15][20][14] = 8'hd6;
frames[15][20][15] = 8'hb5;
frames[15][20][16] = 8'hd6;
frames[15][20][17] = 8'hd6;
frames[15][20][18] = 8'hd6;
frames[15][20][19] = 8'hd6;
frames[15][20][20] = 8'hb1;
frames[15][20][21] = 8'hd5;
frames[15][20][22] = 8'hb1;
frames[15][20][23] = 8'hb6;
frames[15][20][24] = 8'hb6;
frames[15][20][25] = 8'hb1;
frames[15][20][26] = 8'h44;
frames[15][20][27] = 8'h44;
frames[15][20][28] = 8'h44;
frames[15][20][29] = 8'h44;
frames[15][20][30] = 8'h48;
frames[15][20][31] = 8'h48;
frames[15][20][32] = 8'h48;
frames[15][20][33] = 8'h24;
frames[15][20][34] = 8'h48;
frames[15][20][35] = 8'hb6;
frames[15][20][36] = 8'hd6;
frames[15][20][37] = 8'hd6;
frames[15][20][38] = 8'hd6;
frames[15][20][39] = 8'hd6;
frames[15][21][0] = 8'h24;
frames[15][21][1] = 8'h49;
frames[15][21][2] = 8'h44;
frames[15][21][3] = 8'h49;
frames[15][21][4] = 8'hb1;
frames[15][21][5] = 8'hd6;
frames[15][21][6] = 8'hd5;
frames[15][21][7] = 8'hd6;
frames[15][21][8] = 8'hd5;
frames[15][21][9] = 8'hd5;
frames[15][21][10] = 8'hb5;
frames[15][21][11] = 8'hd5;
frames[15][21][12] = 8'hb1;
frames[15][21][13] = 8'hb1;
frames[15][21][14] = 8'hb1;
frames[15][21][15] = 8'h8d;
frames[15][21][16] = 8'hb1;
frames[15][21][17] = 8'hd6;
frames[15][21][18] = 8'hd6;
frames[15][21][19] = 8'hd6;
frames[15][21][20] = 8'hd6;
frames[15][21][21] = 8'hd6;
frames[15][21][22] = 8'hd6;
frames[15][21][23] = 8'hd6;
frames[15][21][24] = 8'hb1;
frames[15][21][25] = 8'h68;
frames[15][21][26] = 8'h44;
frames[15][21][27] = 8'h44;
frames[15][21][28] = 8'h44;
frames[15][21][29] = 8'h44;
frames[15][21][30] = 8'h44;
frames[15][21][31] = 8'h48;
frames[15][21][32] = 8'h48;
frames[15][21][33] = 8'h44;
frames[15][21][34] = 8'h48;
frames[15][21][35] = 8'h91;
frames[15][21][36] = 8'hb2;
frames[15][21][37] = 8'hb2;
frames[15][21][38] = 8'hb2;
frames[15][21][39] = 8'hb6;
frames[15][22][0] = 8'h24;
frames[15][22][1] = 8'h49;
frames[15][22][2] = 8'h48;
frames[15][22][3] = 8'h44;
frames[15][22][4] = 8'h44;
frames[15][22][5] = 8'h69;
frames[15][22][6] = 8'h91;
frames[15][22][7] = 8'hd6;
frames[15][22][8] = 8'hda;
frames[15][22][9] = 8'hd6;
frames[15][22][10] = 8'hb5;
frames[15][22][11] = 8'hd5;
frames[15][22][12] = 8'had;
frames[15][22][13] = 8'had;
frames[15][22][14] = 8'hb1;
frames[15][22][15] = 8'hb1;
frames[15][22][16] = 8'hb5;
frames[15][22][17] = 8'hd6;
frames[15][22][18] = 8'hd6;
frames[15][22][19] = 8'hd6;
frames[15][22][20] = 8'hb5;
frames[15][22][21] = 8'hb1;
frames[15][22][22] = 8'hb1;
frames[15][22][23] = 8'h8d;
frames[15][22][24] = 8'h44;
frames[15][22][25] = 8'h24;
frames[15][22][26] = 8'h44;
frames[15][22][27] = 8'h44;
frames[15][22][28] = 8'h44;
frames[15][22][29] = 8'h48;
frames[15][22][30] = 8'h48;
frames[15][22][31] = 8'h48;
frames[15][22][32] = 8'h48;
frames[15][22][33] = 8'h48;
frames[15][22][34] = 8'h69;
frames[15][22][35] = 8'h6d;
frames[15][22][36] = 8'h8d;
frames[15][22][37] = 8'h8d;
frames[15][22][38] = 8'hb1;
frames[15][22][39] = 8'hb1;
frames[15][23][0] = 8'h49;
frames[15][23][1] = 8'h69;
frames[15][23][2] = 8'h48;
frames[15][23][3] = 8'h48;
frames[15][23][4] = 8'h24;
frames[15][23][5] = 8'h20;
frames[15][23][6] = 8'h20;
frames[15][23][7] = 8'h44;
frames[15][23][8] = 8'h48;
frames[15][23][9] = 8'h6d;
frames[15][23][10] = 8'h8d;
frames[15][23][11] = 8'h91;
frames[15][23][12] = 8'h8d;
frames[15][23][13] = 8'h8d;
frames[15][23][14] = 8'h8d;
frames[15][23][15] = 8'h6c;
frames[15][23][16] = 8'h6d;
frames[15][23][17] = 8'h6d;
frames[15][23][18] = 8'h68;
frames[15][23][19] = 8'h68;
frames[15][23][20] = 8'h48;
frames[15][23][21] = 8'h48;
frames[15][23][22] = 8'h48;
frames[15][23][23] = 8'h44;
frames[15][23][24] = 8'h44;
frames[15][23][25] = 8'h49;
frames[15][23][26] = 8'h49;
frames[15][23][27] = 8'h69;
frames[15][23][28] = 8'h49;
frames[15][23][29] = 8'h49;
frames[15][23][30] = 8'h48;
frames[15][23][31] = 8'h48;
frames[15][23][32] = 8'h44;
frames[15][23][33] = 8'h44;
frames[15][23][34] = 8'h69;
frames[15][23][35] = 8'h6d;
frames[15][23][36] = 8'h8d;
frames[15][23][37] = 8'h8d;
frames[15][23][38] = 8'h8d;
frames[15][23][39] = 8'hb1;
frames[15][24][0] = 8'h48;
frames[15][24][1] = 8'h49;
frames[15][24][2] = 8'h49;
frames[15][24][3] = 8'h48;
frames[15][24][4] = 8'h44;
frames[15][24][5] = 8'h24;
frames[15][24][6] = 8'h24;
frames[15][24][7] = 8'h24;
frames[15][24][8] = 8'h24;
frames[15][24][9] = 8'h24;
frames[15][24][10] = 8'h24;
frames[15][24][11] = 8'h44;
frames[15][24][12] = 8'h44;
frames[15][24][13] = 8'h24;
frames[15][24][14] = 8'h24;
frames[15][24][15] = 8'h24;
frames[15][24][16] = 8'h24;
frames[15][24][17] = 8'h44;
frames[15][24][18] = 8'h44;
frames[15][24][19] = 8'h44;
frames[15][24][20] = 8'h44;
frames[15][24][21] = 8'h44;
frames[15][24][22] = 8'h44;
frames[15][24][23] = 8'h48;
frames[15][24][24] = 8'h48;
frames[15][24][25] = 8'h44;
frames[15][24][26] = 8'h44;
frames[15][24][27] = 8'h44;
frames[15][24][28] = 8'h44;
frames[15][24][29] = 8'h44;
frames[15][24][30] = 8'h24;
frames[15][24][31] = 8'h24;
frames[15][24][32] = 8'h24;
frames[15][24][33] = 8'h24;
frames[15][24][34] = 8'h68;
frames[15][24][35] = 8'h69;
frames[15][24][36] = 8'h69;
frames[15][24][37] = 8'h8d;
frames[15][24][38] = 8'h8d;
frames[15][24][39] = 8'h8d;
frames[15][25][0] = 8'h24;
frames[15][25][1] = 8'h44;
frames[15][25][2] = 8'h44;
frames[15][25][3] = 8'h44;
frames[15][25][4] = 8'h24;
frames[15][25][5] = 8'h24;
frames[15][25][6] = 8'h44;
frames[15][25][7] = 8'h44;
frames[15][25][8] = 8'h24;
frames[15][25][9] = 8'h24;
frames[15][25][10] = 8'h24;
frames[15][25][11] = 8'h24;
frames[15][25][12] = 8'h24;
frames[15][25][13] = 8'h24;
frames[15][25][14] = 8'h24;
frames[15][25][15] = 8'h24;
frames[15][25][16] = 8'h24;
frames[15][25][17] = 8'h24;
frames[15][25][18] = 8'h24;
frames[15][25][19] = 8'h24;
frames[15][25][20] = 8'h24;
frames[15][25][21] = 8'h24;
frames[15][25][22] = 8'h24;
frames[15][25][23] = 8'h24;
frames[15][25][24] = 8'h24;
frames[15][25][25] = 8'h24;
frames[15][25][26] = 8'h24;
frames[15][25][27] = 8'h24;
frames[15][25][28] = 8'h24;
frames[15][25][29] = 8'h24;
frames[15][25][30] = 8'h24;
frames[15][25][31] = 8'h24;
frames[15][25][32] = 8'h44;
frames[15][25][33] = 8'h44;
frames[15][25][34] = 8'h68;
frames[15][25][35] = 8'h68;
frames[15][25][36] = 8'h69;
frames[15][25][37] = 8'h69;
frames[15][25][38] = 8'h8d;
frames[15][25][39] = 8'h8d;
frames[15][26][0] = 8'h24;
frames[15][26][1] = 8'h24;
frames[15][26][2] = 8'h24;
frames[15][26][3] = 8'h24;
frames[15][26][4] = 8'h24;
frames[15][26][5] = 8'h24;
frames[15][26][6] = 8'h24;
frames[15][26][7] = 8'h24;
frames[15][26][8] = 8'h24;
frames[15][26][9] = 8'h24;
frames[15][26][10] = 8'h24;
frames[15][26][11] = 8'h24;
frames[15][26][12] = 8'h24;
frames[15][26][13] = 8'h24;
frames[15][26][14] = 8'h44;
frames[15][26][15] = 8'h44;
frames[15][26][16] = 8'h44;
frames[15][26][17] = 8'h44;
frames[15][26][18] = 8'h44;
frames[15][26][19] = 8'h44;
frames[15][26][20] = 8'h44;
frames[15][26][21] = 8'h44;
frames[15][26][22] = 8'h44;
frames[15][26][23] = 8'h44;
frames[15][26][24] = 8'h44;
frames[15][26][25] = 8'h44;
frames[15][26][26] = 8'h44;
frames[15][26][27] = 8'h44;
frames[15][26][28] = 8'h44;
frames[15][26][29] = 8'h44;
frames[15][26][30] = 8'h44;
frames[15][26][31] = 8'h44;
frames[15][26][32] = 8'h64;
frames[15][26][33] = 8'h68;
frames[15][26][34] = 8'h68;
frames[15][26][35] = 8'h88;
frames[15][26][36] = 8'h88;
frames[15][26][37] = 8'h88;
frames[15][26][38] = 8'h8d;
frames[15][26][39] = 8'h8d;
frames[15][27][0] = 8'h44;
frames[15][27][1] = 8'h44;
frames[15][27][2] = 8'h44;
frames[15][27][3] = 8'h44;
frames[15][27][4] = 8'h44;
frames[15][27][5] = 8'h44;
frames[15][27][6] = 8'h44;
frames[15][27][7] = 8'h44;
frames[15][27][8] = 8'h44;
frames[15][27][9] = 8'h44;
frames[15][27][10] = 8'h44;
frames[15][27][11] = 8'h44;
frames[15][27][12] = 8'h44;
frames[15][27][13] = 8'h44;
frames[15][27][14] = 8'h44;
frames[15][27][15] = 8'h44;
frames[15][27][16] = 8'h44;
frames[15][27][17] = 8'h44;
frames[15][27][18] = 8'h44;
frames[15][27][19] = 8'h44;
frames[15][27][20] = 8'h44;
frames[15][27][21] = 8'h44;
frames[15][27][22] = 8'h64;
frames[15][27][23] = 8'h64;
frames[15][27][24] = 8'h64;
frames[15][27][25] = 8'h64;
frames[15][27][26] = 8'h64;
frames[15][27][27] = 8'h64;
frames[15][27][28] = 8'h64;
frames[15][27][29] = 8'h68;
frames[15][27][30] = 8'h68;
frames[15][27][31] = 8'h68;
frames[15][27][32] = 8'h88;
frames[15][27][33] = 8'h88;
frames[15][27][34] = 8'h88;
frames[15][27][35] = 8'h8c;
frames[15][27][36] = 8'h8c;
frames[15][27][37] = 8'h88;
frames[15][27][38] = 8'h8c;
frames[15][27][39] = 8'h8d;
frames[15][28][0] = 8'h68;
frames[15][28][1] = 8'h68;
frames[15][28][2] = 8'h68;
frames[15][28][3] = 8'h68;
frames[15][28][4] = 8'h68;
frames[15][28][5] = 8'h68;
frames[15][28][6] = 8'h68;
frames[15][28][7] = 8'h68;
frames[15][28][8] = 8'h68;
frames[15][28][9] = 8'h68;
frames[15][28][10] = 8'h68;
frames[15][28][11] = 8'h68;
frames[15][28][12] = 8'h68;
frames[15][28][13] = 8'h68;
frames[15][28][14] = 8'h88;
frames[15][28][15] = 8'h88;
frames[15][28][16] = 8'h88;
frames[15][28][17] = 8'h88;
frames[15][28][18] = 8'h68;
frames[15][28][19] = 8'h68;
frames[15][28][20] = 8'h68;
frames[15][28][21] = 8'h88;
frames[15][28][22] = 8'h88;
frames[15][28][23] = 8'h88;
frames[15][28][24] = 8'h88;
frames[15][28][25] = 8'h68;
frames[15][28][26] = 8'h68;
frames[15][28][27] = 8'h68;
frames[15][28][28] = 8'h68;
frames[15][28][29] = 8'h68;
frames[15][28][30] = 8'h88;
frames[15][28][31] = 8'h88;
frames[15][28][32] = 8'h88;
frames[15][28][33] = 8'h88;
frames[15][28][34] = 8'h8c;
frames[15][28][35] = 8'h8c;
frames[15][28][36] = 8'h8c;
frames[15][28][37] = 8'h88;
frames[15][28][38] = 8'h88;
frames[15][28][39] = 8'h8c;
frames[15][29][0] = 8'h88;
frames[15][29][1] = 8'h88;
frames[15][29][2] = 8'h88;
frames[15][29][3] = 8'h88;
frames[15][29][4] = 8'h88;
frames[15][29][5] = 8'h88;
frames[15][29][6] = 8'h88;
frames[15][29][7] = 8'h88;
frames[15][29][8] = 8'h88;
frames[15][29][9] = 8'h88;
frames[15][29][10] = 8'h88;
frames[15][29][11] = 8'h88;
frames[15][29][12] = 8'h88;
frames[15][29][13] = 8'h8c;
frames[15][29][14] = 8'h8c;
frames[15][29][15] = 8'h8c;
frames[15][29][16] = 8'h8c;
frames[15][29][17] = 8'h88;
frames[15][29][18] = 8'h88;
frames[15][29][19] = 8'h88;
frames[15][29][20] = 8'h88;
frames[15][29][21] = 8'h88;
frames[15][29][22] = 8'h88;
frames[15][29][23] = 8'h88;
frames[15][29][24] = 8'h88;
frames[15][29][25] = 8'h88;
frames[15][29][26] = 8'h88;
frames[15][29][27] = 8'h88;
frames[15][29][28] = 8'h88;
frames[15][29][29] = 8'h88;
frames[15][29][30] = 8'h88;
frames[15][29][31] = 8'h8c;
frames[15][29][32] = 8'h8c;
frames[15][29][33] = 8'h8c;
frames[15][29][34] = 8'h8c;
frames[15][29][35] = 8'hac;
frames[15][29][36] = 8'h8c;
frames[15][29][37] = 8'h88;
frames[15][29][38] = 8'h88;
frames[15][29][39] = 8'h8c;
frames[16][0][0] = 8'had;
frames[16][0][1] = 8'h89;
frames[16][0][2] = 8'h69;
frames[16][0][3] = 8'h20;
frames[16][0][4] = 8'h00;
frames[16][0][5] = 8'h00;
frames[16][0][6] = 8'h00;
frames[16][0][7] = 8'h00;
frames[16][0][8] = 8'h00;
frames[16][0][9] = 8'h00;
frames[16][0][10] = 8'h00;
frames[16][0][11] = 8'h00;
frames[16][0][12] = 8'h00;
frames[16][0][13] = 8'h00;
frames[16][0][14] = 8'h00;
frames[16][0][15] = 8'h00;
frames[16][0][16] = 8'h00;
frames[16][0][17] = 8'h00;
frames[16][0][18] = 8'h00;
frames[16][0][19] = 8'h00;
frames[16][0][20] = 8'h00;
frames[16][0][21] = 8'h00;
frames[16][0][22] = 8'h00;
frames[16][0][23] = 8'h00;
frames[16][0][24] = 8'h00;
frames[16][0][25] = 8'h00;
frames[16][0][26] = 8'h00;
frames[16][0][27] = 8'h24;
frames[16][0][28] = 8'had;
frames[16][0][29] = 8'had;
frames[16][0][30] = 8'ha9;
frames[16][0][31] = 8'ha9;
frames[16][0][32] = 8'h89;
frames[16][0][33] = 8'had;
frames[16][0][34] = 8'h69;
frames[16][0][35] = 8'h69;
frames[16][0][36] = 8'hda;
frames[16][0][37] = 8'hfb;
frames[16][0][38] = 8'hdb;
frames[16][0][39] = 8'hda;
frames[16][1][0] = 8'h89;
frames[16][1][1] = 8'h89;
frames[16][1][2] = 8'h8d;
frames[16][1][3] = 8'h44;
frames[16][1][4] = 8'h00;
frames[16][1][5] = 8'h00;
frames[16][1][6] = 8'h00;
frames[16][1][7] = 8'h00;
frames[16][1][8] = 8'h00;
frames[16][1][9] = 8'h00;
frames[16][1][10] = 8'h00;
frames[16][1][11] = 8'h00;
frames[16][1][12] = 8'h00;
frames[16][1][13] = 8'h00;
frames[16][1][14] = 8'h00;
frames[16][1][15] = 8'h00;
frames[16][1][16] = 8'h00;
frames[16][1][17] = 8'h00;
frames[16][1][18] = 8'h00;
frames[16][1][19] = 8'h00;
frames[16][1][20] = 8'h00;
frames[16][1][21] = 8'h00;
frames[16][1][22] = 8'h00;
frames[16][1][23] = 8'h00;
frames[16][1][24] = 8'h00;
frames[16][1][25] = 8'h00;
frames[16][1][26] = 8'h00;
frames[16][1][27] = 8'h69;
frames[16][1][28] = 8'had;
frames[16][1][29] = 8'ha9;
frames[16][1][30] = 8'h89;
frames[16][1][31] = 8'ha9;
frames[16][1][32] = 8'h89;
frames[16][1][33] = 8'h8d;
frames[16][1][34] = 8'h44;
frames[16][1][35] = 8'h44;
frames[16][1][36] = 8'hdb;
frames[16][1][37] = 8'hfb;
frames[16][1][38] = 8'hdb;
frames[16][1][39] = 8'hdb;
frames[16][2][0] = 8'h89;
frames[16][2][1] = 8'h89;
frames[16][2][2] = 8'h89;
frames[16][2][3] = 8'h88;
frames[16][2][4] = 8'h20;
frames[16][2][5] = 8'h00;
frames[16][2][6] = 8'h00;
frames[16][2][7] = 8'h00;
frames[16][2][8] = 8'h00;
frames[16][2][9] = 8'h00;
frames[16][2][10] = 8'h00;
frames[16][2][11] = 8'h00;
frames[16][2][12] = 8'h00;
frames[16][2][13] = 8'h00;
frames[16][2][14] = 8'h00;
frames[16][2][15] = 8'h00;
frames[16][2][16] = 8'h00;
frames[16][2][17] = 8'h00;
frames[16][2][18] = 8'h00;
frames[16][2][19] = 8'h00;
frames[16][2][20] = 8'h00;
frames[16][2][21] = 8'h00;
frames[16][2][22] = 8'h00;
frames[16][2][23] = 8'h00;
frames[16][2][24] = 8'h00;
frames[16][2][25] = 8'h00;
frames[16][2][26] = 8'h20;
frames[16][2][27] = 8'h8d;
frames[16][2][28] = 8'had;
frames[16][2][29] = 8'had;
frames[16][2][30] = 8'ha9;
frames[16][2][31] = 8'ha9;
frames[16][2][32] = 8'h8d;
frames[16][2][33] = 8'h89;
frames[16][2][34] = 8'h20;
frames[16][2][35] = 8'h24;
frames[16][2][36] = 8'hdb;
frames[16][2][37] = 8'hdb;
frames[16][2][38] = 8'h49;
frames[16][2][39] = 8'hbb;
frames[16][3][0] = 8'h89;
frames[16][3][1] = 8'h89;
frames[16][3][2] = 8'h89;
frames[16][3][3] = 8'h89;
frames[16][3][4] = 8'h44;
frames[16][3][5] = 8'h00;
frames[16][3][6] = 8'h00;
frames[16][3][7] = 8'h00;
frames[16][3][8] = 8'h00;
frames[16][3][9] = 8'h00;
frames[16][3][10] = 8'h00;
frames[16][3][11] = 8'h00;
frames[16][3][12] = 8'h00;
frames[16][3][13] = 8'h00;
frames[16][3][14] = 8'h00;
frames[16][3][15] = 8'h00;
frames[16][3][16] = 8'h00;
frames[16][3][17] = 8'h00;
frames[16][3][18] = 8'h00;
frames[16][3][19] = 8'h00;
frames[16][3][20] = 8'h00;
frames[16][3][21] = 8'h00;
frames[16][3][22] = 8'h00;
frames[16][3][23] = 8'h00;
frames[16][3][24] = 8'h00;
frames[16][3][25] = 8'h00;
frames[16][3][26] = 8'h44;
frames[16][3][27] = 8'h8d;
frames[16][3][28] = 8'had;
frames[16][3][29] = 8'ha9;
frames[16][3][30] = 8'ha9;
frames[16][3][31] = 8'ha9;
frames[16][3][32] = 8'ha9;
frames[16][3][33] = 8'had;
frames[16][3][34] = 8'h24;
frames[16][3][35] = 8'h20;
frames[16][3][36] = 8'hdb;
frames[16][3][37] = 8'hdb;
frames[16][3][38] = 8'h49;
frames[16][3][39] = 8'hb7;
frames[16][4][0] = 8'ha9;
frames[16][4][1] = 8'ha9;
frames[16][4][2] = 8'h89;
frames[16][4][3] = 8'h89;
frames[16][4][4] = 8'h69;
frames[16][4][5] = 8'h20;
frames[16][4][6] = 8'h00;
frames[16][4][7] = 8'h00;
frames[16][4][8] = 8'h00;
frames[16][4][9] = 8'h00;
frames[16][4][10] = 8'h00;
frames[16][4][11] = 8'h00;
frames[16][4][12] = 8'h00;
frames[16][4][13] = 8'h00;
frames[16][4][14] = 8'h00;
frames[16][4][15] = 8'h00;
frames[16][4][16] = 8'h00;
frames[16][4][17] = 8'h00;
frames[16][4][18] = 8'h00;
frames[16][4][19] = 8'h00;
frames[16][4][20] = 8'h00;
frames[16][4][21] = 8'h00;
frames[16][4][22] = 8'h00;
frames[16][4][23] = 8'h00;
frames[16][4][24] = 8'h00;
frames[16][4][25] = 8'h00;
frames[16][4][26] = 8'h44;
frames[16][4][27] = 8'h8d;
frames[16][4][28] = 8'ha9;
frames[16][4][29] = 8'ha9;
frames[16][4][30] = 8'h89;
frames[16][4][31] = 8'ha9;
frames[16][4][32] = 8'had;
frames[16][4][33] = 8'had;
frames[16][4][34] = 8'h69;
frames[16][4][35] = 8'h00;
frames[16][4][36] = 8'hb6;
frames[16][4][37] = 8'hdb;
frames[16][4][38] = 8'h6e;
frames[16][4][39] = 8'hdb;
frames[16][5][0] = 8'had;
frames[16][5][1] = 8'had;
frames[16][5][2] = 8'h89;
frames[16][5][3] = 8'h89;
frames[16][5][4] = 8'h69;
frames[16][5][5] = 8'h20;
frames[16][5][6] = 8'h00;
frames[16][5][7] = 8'h00;
frames[16][5][8] = 8'h00;
frames[16][5][9] = 8'h00;
frames[16][5][10] = 8'h00;
frames[16][5][11] = 8'h00;
frames[16][5][12] = 8'h00;
frames[16][5][13] = 8'h00;
frames[16][5][14] = 8'h00;
frames[16][5][15] = 8'h00;
frames[16][5][16] = 8'h00;
frames[16][5][17] = 8'h00;
frames[16][5][18] = 8'h00;
frames[16][5][19] = 8'h00;
frames[16][5][20] = 8'h00;
frames[16][5][21] = 8'h00;
frames[16][5][22] = 8'h00;
frames[16][5][23] = 8'h00;
frames[16][5][24] = 8'h00;
frames[16][5][25] = 8'h00;
frames[16][5][26] = 8'h68;
frames[16][5][27] = 8'h8d;
frames[16][5][28] = 8'h89;
frames[16][5][29] = 8'h88;
frames[16][5][30] = 8'h89;
frames[16][5][31] = 8'had;
frames[16][5][32] = 8'had;
frames[16][5][33] = 8'had;
frames[16][5][34] = 8'h8d;
frames[16][5][35] = 8'h20;
frames[16][5][36] = 8'h6d;
frames[16][5][37] = 8'hfb;
frames[16][5][38] = 8'hdb;
frames[16][5][39] = 8'hdb;
frames[16][6][0] = 8'had;
frames[16][6][1] = 8'had;
frames[16][6][2] = 8'h89;
frames[16][6][3] = 8'h89;
frames[16][6][4] = 8'h69;
frames[16][6][5] = 8'h20;
frames[16][6][6] = 8'h00;
frames[16][6][7] = 8'h00;
frames[16][6][8] = 8'h00;
frames[16][6][9] = 8'h00;
frames[16][6][10] = 8'h00;
frames[16][6][11] = 8'h00;
frames[16][6][12] = 8'h00;
frames[16][6][13] = 8'h00;
frames[16][6][14] = 8'h00;
frames[16][6][15] = 8'h00;
frames[16][6][16] = 8'h00;
frames[16][6][17] = 8'h00;
frames[16][6][18] = 8'h00;
frames[16][6][19] = 8'h00;
frames[16][6][20] = 8'h00;
frames[16][6][21] = 8'h00;
frames[16][6][22] = 8'h00;
frames[16][6][23] = 8'h00;
frames[16][6][24] = 8'h00;
frames[16][6][25] = 8'h00;
frames[16][6][26] = 8'h89;
frames[16][6][27] = 8'ha9;
frames[16][6][28] = 8'h89;
frames[16][6][29] = 8'h64;
frames[16][6][30] = 8'h89;
frames[16][6][31] = 8'had;
frames[16][6][32] = 8'had;
frames[16][6][33] = 8'had;
frames[16][6][34] = 8'h8d;
frames[16][6][35] = 8'h44;
frames[16][6][36] = 8'h48;
frames[16][6][37] = 8'hda;
frames[16][6][38] = 8'hda;
frames[16][6][39] = 8'hda;
frames[16][7][0] = 8'h89;
frames[16][7][1] = 8'h89;
frames[16][7][2] = 8'h89;
frames[16][7][3] = 8'h89;
frames[16][7][4] = 8'h69;
frames[16][7][5] = 8'h20;
frames[16][7][6] = 8'h00;
frames[16][7][7] = 8'h00;
frames[16][7][8] = 8'h00;
frames[16][7][9] = 8'h00;
frames[16][7][10] = 8'h00;
frames[16][7][11] = 8'h00;
frames[16][7][12] = 8'h00;
frames[16][7][13] = 8'h00;
frames[16][7][14] = 8'h00;
frames[16][7][15] = 8'h00;
frames[16][7][16] = 8'h00;
frames[16][7][17] = 8'h00;
frames[16][7][18] = 8'h00;
frames[16][7][19] = 8'h00;
frames[16][7][20] = 8'h00;
frames[16][7][21] = 8'h00;
frames[16][7][22] = 8'h00;
frames[16][7][23] = 8'h00;
frames[16][7][24] = 8'h00;
frames[16][7][25] = 8'h20;
frames[16][7][26] = 8'h89;
frames[16][7][27] = 8'h89;
frames[16][7][28] = 8'h64;
frames[16][7][29] = 8'h40;
frames[16][7][30] = 8'had;
frames[16][7][31] = 8'had;
frames[16][7][32] = 8'had;
frames[16][7][33] = 8'had;
frames[16][7][34] = 8'had;
frames[16][7][35] = 8'h68;
frames[16][7][36] = 8'h44;
frames[16][7][37] = 8'hdb;
frames[16][7][38] = 8'hdb;
frames[16][7][39] = 8'hdb;
frames[16][8][0] = 8'h84;
frames[16][8][1] = 8'h88;
frames[16][8][2] = 8'h88;
frames[16][8][3] = 8'h89;
frames[16][8][4] = 8'h89;
frames[16][8][5] = 8'h40;
frames[16][8][6] = 8'h00;
frames[16][8][7] = 8'h00;
frames[16][8][8] = 8'h00;
frames[16][8][9] = 8'h00;
frames[16][8][10] = 8'h00;
frames[16][8][11] = 8'h00;
frames[16][8][12] = 8'h00;
frames[16][8][13] = 8'h00;
frames[16][8][14] = 8'h00;
frames[16][8][15] = 8'h00;
frames[16][8][16] = 8'h00;
frames[16][8][17] = 8'h00;
frames[16][8][18] = 8'h00;
frames[16][8][19] = 8'h00;
frames[16][8][20] = 8'h00;
frames[16][8][21] = 8'h00;
frames[16][8][22] = 8'h00;
frames[16][8][23] = 8'h00;
frames[16][8][24] = 8'h00;
frames[16][8][25] = 8'h44;
frames[16][8][26] = 8'had;
frames[16][8][27] = 8'h89;
frames[16][8][28] = 8'h40;
frames[16][8][29] = 8'h64;
frames[16][8][30] = 8'had;
frames[16][8][31] = 8'had;
frames[16][8][32] = 8'had;
frames[16][8][33] = 8'had;
frames[16][8][34] = 8'had;
frames[16][8][35] = 8'h68;
frames[16][8][36] = 8'h24;
frames[16][8][37] = 8'hdb;
frames[16][8][38] = 8'hda;
frames[16][8][39] = 8'hda;
frames[16][9][0] = 8'h64;
frames[16][9][1] = 8'h64;
frames[16][9][2] = 8'h64;
frames[16][9][3] = 8'h88;
frames[16][9][4] = 8'h89;
frames[16][9][5] = 8'h44;
frames[16][9][6] = 8'h00;
frames[16][9][7] = 8'h20;
frames[16][9][8] = 8'h44;
frames[16][9][9] = 8'h69;
frames[16][9][10] = 8'h69;
frames[16][9][11] = 8'h6d;
frames[16][9][12] = 8'h8d;
frames[16][9][13] = 8'h8d;
frames[16][9][14] = 8'h8d;
frames[16][9][15] = 8'h8d;
frames[16][9][16] = 8'h69;
frames[16][9][17] = 8'h68;
frames[16][9][18] = 8'h69;
frames[16][9][19] = 8'h48;
frames[16][9][20] = 8'h24;
frames[16][9][21] = 8'h24;
frames[16][9][22] = 8'h24;
frames[16][9][23] = 8'h24;
frames[16][9][24] = 8'h44;
frames[16][9][25] = 8'h69;
frames[16][9][26] = 8'h89;
frames[16][9][27] = 8'h88;
frames[16][9][28] = 8'h64;
frames[16][9][29] = 8'h8d;
frames[16][9][30] = 8'had;
frames[16][9][31] = 8'had;
frames[16][9][32] = 8'had;
frames[16][9][33] = 8'had;
frames[16][9][34] = 8'h8d;
frames[16][9][35] = 8'h44;
frames[16][9][36] = 8'h6d;
frames[16][9][37] = 8'hfb;
frames[16][9][38] = 8'hdb;
frames[16][9][39] = 8'hda;
frames[16][10][0] = 8'h68;
frames[16][10][1] = 8'h44;
frames[16][10][2] = 8'h20;
frames[16][10][3] = 8'h44;
frames[16][10][4] = 8'h89;
frames[16][10][5] = 8'h64;
frames[16][10][6] = 8'h48;
frames[16][10][7] = 8'h8d;
frames[16][10][8] = 8'hb1;
frames[16][10][9] = 8'hb1;
frames[16][10][10] = 8'hb1;
frames[16][10][11] = 8'hb1;
frames[16][10][12] = 8'hd1;
frames[16][10][13] = 8'hb1;
frames[16][10][14] = 8'hb1;
frames[16][10][15] = 8'hb1;
frames[16][10][16] = 8'hb1;
frames[16][10][17] = 8'hb1;
frames[16][10][18] = 8'hb1;
frames[16][10][19] = 8'hb1;
frames[16][10][20] = 8'h91;
frames[16][10][21] = 8'h8d;
frames[16][10][22] = 8'h6d;
frames[16][10][23] = 8'h6d;
frames[16][10][24] = 8'h89;
frames[16][10][25] = 8'h8d;
frames[16][10][26] = 8'h89;
frames[16][10][27] = 8'h64;
frames[16][10][28] = 8'h89;
frames[16][10][29] = 8'had;
frames[16][10][30] = 8'had;
frames[16][10][31] = 8'had;
frames[16][10][32] = 8'had;
frames[16][10][33] = 8'had;
frames[16][10][34] = 8'h44;
frames[16][10][35] = 8'h69;
frames[16][10][36] = 8'hdb;
frames[16][10][37] = 8'hff;
frames[16][10][38] = 8'hdb;
frames[16][10][39] = 8'hda;
frames[16][11][0] = 8'h89;
frames[16][11][1] = 8'h64;
frames[16][11][2] = 8'h20;
frames[16][11][3] = 8'h44;
frames[16][11][4] = 8'h88;
frames[16][11][5] = 8'h89;
frames[16][11][6] = 8'had;
frames[16][11][7] = 8'hb1;
frames[16][11][8] = 8'hb1;
frames[16][11][9] = 8'hb1;
frames[16][11][10] = 8'hb1;
frames[16][11][11] = 8'hb1;
frames[16][11][12] = 8'hb1;
frames[16][11][13] = 8'hb1;
frames[16][11][14] = 8'hb1;
frames[16][11][15] = 8'hb1;
frames[16][11][16] = 8'hb1;
frames[16][11][17] = 8'hb1;
frames[16][11][18] = 8'hb5;
frames[16][11][19] = 8'hb1;
frames[16][11][20] = 8'hb1;
frames[16][11][21] = 8'hb1;
frames[16][11][22] = 8'hb1;
frames[16][11][23] = 8'hb1;
frames[16][11][24] = 8'had;
frames[16][11][25] = 8'h89;
frames[16][11][26] = 8'h84;
frames[16][11][27] = 8'h88;
frames[16][11][28] = 8'had;
frames[16][11][29] = 8'had;
frames[16][11][30] = 8'h89;
frames[16][11][31] = 8'had;
frames[16][11][32] = 8'had;
frames[16][11][33] = 8'h89;
frames[16][11][34] = 8'h24;
frames[16][11][35] = 8'h6d;
frames[16][11][36] = 8'hdb;
frames[16][11][37] = 8'hff;
frames[16][11][38] = 8'hdb;
frames[16][11][39] = 8'hda;
frames[16][12][0] = 8'h89;
frames[16][12][1] = 8'h89;
frames[16][12][2] = 8'h44;
frames[16][12][3] = 8'h40;
frames[16][12][4] = 8'h64;
frames[16][12][5] = 8'h89;
frames[16][12][6] = 8'h8d;
frames[16][12][7] = 8'hb1;
frames[16][12][8] = 8'hb1;
frames[16][12][9] = 8'hb1;
frames[16][12][10] = 8'hb1;
frames[16][12][11] = 8'hb1;
frames[16][12][12] = 8'hb1;
frames[16][12][13] = 8'hb1;
frames[16][12][14] = 8'hb1;
frames[16][12][15] = 8'hb1;
frames[16][12][16] = 8'hb1;
frames[16][12][17] = 8'hb1;
frames[16][12][18] = 8'hb1;
frames[16][12][19] = 8'hb1;
frames[16][12][20] = 8'hb1;
frames[16][12][21] = 8'hb1;
frames[16][12][22] = 8'hb1;
frames[16][12][23] = 8'had;
frames[16][12][24] = 8'h89;
frames[16][12][25] = 8'h89;
frames[16][12][26] = 8'h89;
frames[16][12][27] = 8'had;
frames[16][12][28] = 8'had;
frames[16][12][29] = 8'h89;
frames[16][12][30] = 8'h89;
frames[16][12][31] = 8'had;
frames[16][12][32] = 8'h8d;
frames[16][12][33] = 8'h44;
frames[16][12][34] = 8'h24;
frames[16][12][35] = 8'h91;
frames[16][12][36] = 8'hdb;
frames[16][12][37] = 8'hfb;
frames[16][12][38] = 8'hdb;
frames[16][12][39] = 8'hda;
frames[16][13][0] = 8'h88;
frames[16][13][1] = 8'h89;
frames[16][13][2] = 8'h89;
frames[16][13][3] = 8'h64;
frames[16][13][4] = 8'h64;
frames[16][13][5] = 8'h89;
frames[16][13][6] = 8'h89;
frames[16][13][7] = 8'had;
frames[16][13][8] = 8'hb1;
frames[16][13][9] = 8'hb1;
frames[16][13][10] = 8'hb1;
frames[16][13][11] = 8'hb1;
frames[16][13][12] = 8'hb1;
frames[16][13][13] = 8'hb1;
frames[16][13][14] = 8'hb1;
frames[16][13][15] = 8'hb1;
frames[16][13][16] = 8'hb1;
frames[16][13][17] = 8'hb1;
frames[16][13][18] = 8'hb1;
frames[16][13][19] = 8'hb1;
frames[16][13][20] = 8'h91;
frames[16][13][21] = 8'h91;
frames[16][13][22] = 8'hb1;
frames[16][13][23] = 8'h8d;
frames[16][13][24] = 8'h89;
frames[16][13][25] = 8'had;
frames[16][13][26] = 8'had;
frames[16][13][27] = 8'had;
frames[16][13][28] = 8'had;
frames[16][13][29] = 8'had;
frames[16][13][30] = 8'had;
frames[16][13][31] = 8'had;
frames[16][13][32] = 8'h48;
frames[16][13][33] = 8'h24;
frames[16][13][34] = 8'h44;
frames[16][13][35] = 8'hb2;
frames[16][13][36] = 8'hdb;
frames[16][13][37] = 8'hdb;
frames[16][13][38] = 8'hdb;
frames[16][13][39] = 8'hda;
frames[16][14][0] = 8'h88;
frames[16][14][1] = 8'h88;
frames[16][14][2] = 8'h89;
frames[16][14][3] = 8'h89;
frames[16][14][4] = 8'h89;
frames[16][14][5] = 8'h88;
frames[16][14][6] = 8'h8d;
frames[16][14][7] = 8'h8d;
frames[16][14][8] = 8'hb1;
frames[16][14][9] = 8'hb1;
frames[16][14][10] = 8'hb1;
frames[16][14][11] = 8'hb1;
frames[16][14][12] = 8'hb1;
frames[16][14][13] = 8'hb1;
frames[16][14][14] = 8'hb1;
frames[16][14][15] = 8'hb1;
frames[16][14][16] = 8'hb1;
frames[16][14][17] = 8'hb1;
frames[16][14][18] = 8'hb1;
frames[16][14][19] = 8'hb1;
frames[16][14][20] = 8'hb1;
frames[16][14][21] = 8'hb1;
frames[16][14][22] = 8'hb1;
frames[16][14][23] = 8'h8d;
frames[16][14][24] = 8'had;
frames[16][14][25] = 8'had;
frames[16][14][26] = 8'ha9;
frames[16][14][27] = 8'ha9;
frames[16][14][28] = 8'had;
frames[16][14][29] = 8'had;
frames[16][14][30] = 8'h89;
frames[16][14][31] = 8'h64;
frames[16][14][32] = 8'h24;
frames[16][14][33] = 8'h44;
frames[16][14][34] = 8'h49;
frames[16][14][35] = 8'hb6;
frames[16][14][36] = 8'hdb;
frames[16][14][37] = 8'hdb;
frames[16][14][38] = 8'hdb;
frames[16][14][39] = 8'hda;
frames[16][15][0] = 8'had;
frames[16][15][1] = 8'ha9;
frames[16][15][2] = 8'h88;
frames[16][15][3] = 8'h88;
frames[16][15][4] = 8'h89;
frames[16][15][5] = 8'h64;
frames[16][15][6] = 8'h68;
frames[16][15][7] = 8'had;
frames[16][15][8] = 8'hb1;
frames[16][15][9] = 8'hb1;
frames[16][15][10] = 8'h91;
frames[16][15][11] = 8'h91;
frames[16][15][12] = 8'hb1;
frames[16][15][13] = 8'hb1;
frames[16][15][14] = 8'hb1;
frames[16][15][15] = 8'hb1;
frames[16][15][16] = 8'hb1;
frames[16][15][17] = 8'hb1;
frames[16][15][18] = 8'hb1;
frames[16][15][19] = 8'hb1;
frames[16][15][20] = 8'hb1;
frames[16][15][21] = 8'hb1;
frames[16][15][22] = 8'hb1;
frames[16][15][23] = 8'hb1;
frames[16][15][24] = 8'h8d;
frames[16][15][25] = 8'h68;
frames[16][15][26] = 8'h64;
frames[16][15][27] = 8'h68;
frames[16][15][28] = 8'h68;
frames[16][15][29] = 8'h64;
frames[16][15][30] = 8'h44;
frames[16][15][31] = 8'h24;
frames[16][15][32] = 8'h24;
frames[16][15][33] = 8'h44;
frames[16][15][34] = 8'h6d;
frames[16][15][35] = 8'hb6;
frames[16][15][36] = 8'hdb;
frames[16][15][37] = 8'hdb;
frames[16][15][38] = 8'hdb;
frames[16][15][39] = 8'hda;
frames[16][16][0] = 8'h89;
frames[16][16][1] = 8'h89;
frames[16][16][2] = 8'h88;
frames[16][16][3] = 8'h88;
frames[16][16][4] = 8'h88;
frames[16][16][5] = 8'h64;
frames[16][16][6] = 8'h68;
frames[16][16][7] = 8'hb1;
frames[16][16][8] = 8'h91;
frames[16][16][9] = 8'h91;
frames[16][16][10] = 8'hb1;
frames[16][16][11] = 8'hb1;
frames[16][16][12] = 8'hb1;
frames[16][16][13] = 8'hb1;
frames[16][16][14] = 8'hb1;
frames[16][16][15] = 8'hb1;
frames[16][16][16] = 8'hb1;
frames[16][16][17] = 8'hb1;
frames[16][16][18] = 8'hb1;
frames[16][16][19] = 8'hb1;
frames[16][16][20] = 8'hb1;
frames[16][16][21] = 8'hd2;
frames[16][16][22] = 8'hb1;
frames[16][16][23] = 8'h48;
frames[16][16][24] = 8'h24;
frames[16][16][25] = 8'h24;
frames[16][16][26] = 8'h24;
frames[16][16][27] = 8'h24;
frames[16][16][28] = 8'h24;
frames[16][16][29] = 8'h20;
frames[16][16][30] = 8'h24;
frames[16][16][31] = 8'h20;
frames[16][16][32] = 8'h20;
frames[16][16][33] = 8'h24;
frames[16][16][34] = 8'h6d;
frames[16][16][35] = 8'hd6;
frames[16][16][36] = 8'hdb;
frames[16][16][37] = 8'hdb;
frames[16][16][38] = 8'hdb;
frames[16][16][39] = 8'hda;
frames[16][17][0] = 8'h69;
frames[16][17][1] = 8'h44;
frames[16][17][2] = 8'h64;
frames[16][17][3] = 8'h68;
frames[16][17][4] = 8'h68;
frames[16][17][5] = 8'h44;
frames[16][17][6] = 8'h68;
frames[16][17][7] = 8'h8d;
frames[16][17][8] = 8'h8d;
frames[16][17][9] = 8'h8d;
frames[16][17][10] = 8'h8d;
frames[16][17][11] = 8'h91;
frames[16][17][12] = 8'hb1;
frames[16][17][13] = 8'hb1;
frames[16][17][14] = 8'hb1;
frames[16][17][15] = 8'hb1;
frames[16][17][16] = 8'hb1;
frames[16][17][17] = 8'hb1;
frames[16][17][18] = 8'hb1;
frames[16][17][19] = 8'hb1;
frames[16][17][20] = 8'hb1;
frames[16][17][21] = 8'h69;
frames[16][17][22] = 8'h44;
frames[16][17][23] = 8'h24;
frames[16][17][24] = 8'h24;
frames[16][17][25] = 8'h24;
frames[16][17][26] = 8'h24;
frames[16][17][27] = 8'h20;
frames[16][17][28] = 8'h20;
frames[16][17][29] = 8'h20;
frames[16][17][30] = 8'h24;
frames[16][17][31] = 8'h20;
frames[16][17][32] = 8'h20;
frames[16][17][33] = 8'h24;
frames[16][17][34] = 8'h6d;
frames[16][17][35] = 8'hd6;
frames[16][17][36] = 8'hfb;
frames[16][17][37] = 8'hdb;
frames[16][17][38] = 8'hdb;
frames[16][17][39] = 8'hda;
frames[16][18][0] = 8'h49;
frames[16][18][1] = 8'h24;
frames[16][18][2] = 8'h69;
frames[16][18][3] = 8'h69;
frames[16][18][4] = 8'h69;
frames[16][18][5] = 8'h49;
frames[16][18][6] = 8'h48;
frames[16][18][7] = 8'h44;
frames[16][18][8] = 8'h68;
frames[16][18][9] = 8'h68;
frames[16][18][10] = 8'h68;
frames[16][18][11] = 8'h8d;
frames[16][18][12] = 8'h91;
frames[16][18][13] = 8'hb1;
frames[16][18][14] = 8'hb1;
frames[16][18][15] = 8'hb1;
frames[16][18][16] = 8'hb1;
frames[16][18][17] = 8'hb1;
frames[16][18][18] = 8'hb1;
frames[16][18][19] = 8'hb1;
frames[16][18][20] = 8'h8d;
frames[16][18][21] = 8'h69;
frames[16][18][22] = 8'h24;
frames[16][18][23] = 8'h24;
frames[16][18][24] = 8'h24;
frames[16][18][25] = 8'h24;
frames[16][18][26] = 8'h24;
frames[16][18][27] = 8'h20;
frames[16][18][28] = 8'h20;
frames[16][18][29] = 8'h20;
frames[16][18][30] = 8'h24;
frames[16][18][31] = 8'h24;
frames[16][18][32] = 8'h24;
frames[16][18][33] = 8'h20;
frames[16][18][34] = 8'h49;
frames[16][18][35] = 8'hd6;
frames[16][18][36] = 8'hfb;
frames[16][18][37] = 8'hdb;
frames[16][18][38] = 8'hdb;
frames[16][18][39] = 8'hd6;
frames[16][19][0] = 8'h48;
frames[16][19][1] = 8'h24;
frames[16][19][2] = 8'h6d;
frames[16][19][3] = 8'h6d;
frames[16][19][4] = 8'h69;
frames[16][19][5] = 8'h69;
frames[16][19][6] = 8'h69;
frames[16][19][7] = 8'h69;
frames[16][19][8] = 8'h68;
frames[16][19][9] = 8'h6d;
frames[16][19][10] = 8'h6c;
frames[16][19][11] = 8'h8d;
frames[16][19][12] = 8'hb1;
frames[16][19][13] = 8'hb1;
frames[16][19][14] = 8'hb1;
frames[16][19][15] = 8'hb1;
frames[16][19][16] = 8'hb1;
frames[16][19][17] = 8'hb1;
frames[16][19][18] = 8'hb5;
frames[16][19][19] = 8'hb5;
frames[16][19][20] = 8'hd6;
frames[16][19][21] = 8'hb1;
frames[16][19][22] = 8'h8d;
frames[16][19][23] = 8'h69;
frames[16][19][24] = 8'h24;
frames[16][19][25] = 8'h24;
frames[16][19][26] = 8'h24;
frames[16][19][27] = 8'h20;
frames[16][19][28] = 8'h20;
frames[16][19][29] = 8'h20;
frames[16][19][30] = 8'h20;
frames[16][19][31] = 8'h24;
frames[16][19][32] = 8'h24;
frames[16][19][33] = 8'h20;
frames[16][19][34] = 8'h24;
frames[16][19][35] = 8'hb6;
frames[16][19][36] = 8'hfb;
frames[16][19][37] = 8'hdb;
frames[16][19][38] = 8'hdb;
frames[16][19][39] = 8'hd6;
frames[16][20][0] = 8'h24;
frames[16][20][1] = 8'h48;
frames[16][20][2] = 8'h6d;
frames[16][20][3] = 8'h6d;
frames[16][20][4] = 8'h69;
frames[16][20][5] = 8'h6d;
frames[16][20][6] = 8'h8d;
frames[16][20][7] = 8'h8d;
frames[16][20][8] = 8'had;
frames[16][20][9] = 8'h88;
frames[16][20][10] = 8'h68;
frames[16][20][11] = 8'hb1;
frames[16][20][12] = 8'hb1;
frames[16][20][13] = 8'hd5;
frames[16][20][14] = 8'hd5;
frames[16][20][15] = 8'hb5;
frames[16][20][16] = 8'hb1;
frames[16][20][17] = 8'hd5;
frames[16][20][18] = 8'hd6;
frames[16][20][19] = 8'hd6;
frames[16][20][20] = 8'hd6;
frames[16][20][21] = 8'hd6;
frames[16][20][22] = 8'hb1;
frames[16][20][23] = 8'hb1;
frames[16][20][24] = 8'h8d;
frames[16][20][25] = 8'h48;
frames[16][20][26] = 8'h24;
frames[16][20][27] = 8'h24;
frames[16][20][28] = 8'h20;
frames[16][20][29] = 8'h20;
frames[16][20][30] = 8'h24;
frames[16][20][31] = 8'h24;
frames[16][20][32] = 8'h44;
frames[16][20][33] = 8'h20;
frames[16][20][34] = 8'h24;
frames[16][20][35] = 8'h92;
frames[16][20][36] = 8'hfb;
frames[16][20][37] = 8'hdb;
frames[16][20][38] = 8'hdb;
frames[16][20][39] = 8'hd6;
frames[16][21][0] = 8'h24;
frames[16][21][1] = 8'h49;
frames[16][21][2] = 8'h6d;
frames[16][21][3] = 8'h6d;
frames[16][21][4] = 8'h6d;
frames[16][21][5] = 8'h91;
frames[16][21][6] = 8'hb1;
frames[16][21][7] = 8'h8d;
frames[16][21][8] = 8'h88;
frames[16][21][9] = 8'had;
frames[16][21][10] = 8'hb1;
frames[16][21][11] = 8'hd6;
frames[16][21][12] = 8'hb1;
frames[16][21][13] = 8'hb1;
frames[16][21][14] = 8'hb5;
frames[16][21][15] = 8'hd6;
frames[16][21][16] = 8'hd6;
frames[16][21][17] = 8'hd5;
frames[16][21][18] = 8'hd6;
frames[16][21][19] = 8'hb1;
frames[16][21][20] = 8'hb1;
frames[16][21][21] = 8'hd5;
frames[16][21][22] = 8'hb5;
frames[16][21][23] = 8'hd6;
frames[16][21][24] = 8'hb1;
frames[16][21][25] = 8'hb1;
frames[16][21][26] = 8'h6d;
frames[16][21][27] = 8'h48;
frames[16][21][28] = 8'h24;
frames[16][21][29] = 8'h20;
frames[16][21][30] = 8'h24;
frames[16][21][31] = 8'h44;
frames[16][21][32] = 8'h44;
frames[16][21][33] = 8'h24;
frames[16][21][34] = 8'h20;
frames[16][21][35] = 8'h6d;
frames[16][21][36] = 8'hfb;
frames[16][21][37] = 8'hdb;
frames[16][21][38] = 8'hdb;
frames[16][21][39] = 8'hd6;
frames[16][22][0] = 8'h24;
frames[16][22][1] = 8'h49;
frames[16][22][2] = 8'h6d;
frames[16][22][3] = 8'h6d;
frames[16][22][4] = 8'h91;
frames[16][22][5] = 8'hb1;
frames[16][22][6] = 8'hb1;
frames[16][22][7] = 8'h8d;
frames[16][22][8] = 8'h68;
frames[16][22][9] = 8'h88;
frames[16][22][10] = 8'hb1;
frames[16][22][11] = 8'hb5;
frames[16][22][12] = 8'hb5;
frames[16][22][13] = 8'hb1;
frames[16][22][14] = 8'hb1;
frames[16][22][15] = 8'hd5;
frames[16][22][16] = 8'hd5;
frames[16][22][17] = 8'hd6;
frames[16][22][18] = 8'hd6;
frames[16][22][19] = 8'hd6;
frames[16][22][20] = 8'hb5;
frames[16][22][21] = 8'hb1;
frames[16][22][22] = 8'hb1;
frames[16][22][23] = 8'hb1;
frames[16][22][24] = 8'hb5;
frames[16][22][25] = 8'hb5;
frames[16][22][26] = 8'h8d;
frames[16][22][27] = 8'h20;
frames[16][22][28] = 8'h24;
frames[16][22][29] = 8'h20;
frames[16][22][30] = 8'h24;
frames[16][22][31] = 8'h44;
frames[16][22][32] = 8'h44;
frames[16][22][33] = 8'h24;
frames[16][22][34] = 8'h20;
frames[16][22][35] = 8'h48;
frames[16][22][36] = 8'hda;
frames[16][22][37] = 8'hdb;
frames[16][22][38] = 8'hda;
frames[16][22][39] = 8'hd6;
frames[16][23][0] = 8'h24;
frames[16][23][1] = 8'h6d;
frames[16][23][2] = 8'h6d;
frames[16][23][3] = 8'h6d;
frames[16][23][4] = 8'h8d;
frames[16][23][5] = 8'hb2;
frames[16][23][6] = 8'hb1;
frames[16][23][7] = 8'hb1;
frames[16][23][8] = 8'hb1;
frames[16][23][9] = 8'hb1;
frames[16][23][10] = 8'hb1;
frames[16][23][11] = 8'hb1;
frames[16][23][12] = 8'hb1;
frames[16][23][13] = 8'hb1;
frames[16][23][14] = 8'had;
frames[16][23][15] = 8'had;
frames[16][23][16] = 8'h8d;
frames[16][23][17] = 8'hd5;
frames[16][23][18] = 8'hd6;
frames[16][23][19] = 8'hd6;
frames[16][23][20] = 8'hd6;
frames[16][23][21] = 8'hb5;
frames[16][23][22] = 8'hd6;
frames[16][23][23] = 8'hd6;
frames[16][23][24] = 8'hb6;
frames[16][23][25] = 8'hb1;
frames[16][23][26] = 8'h48;
frames[16][23][27] = 8'h20;
frames[16][23][28] = 8'h24;
frames[16][23][29] = 8'h20;
frames[16][23][30] = 8'h24;
frames[16][23][31] = 8'h44;
frames[16][23][32] = 8'h44;
frames[16][23][33] = 8'h44;
frames[16][23][34] = 8'h20;
frames[16][23][35] = 8'h44;
frames[16][23][36] = 8'hb6;
frames[16][23][37] = 8'hda;
frames[16][23][38] = 8'hd6;
frames[16][23][39] = 8'hd6;
frames[16][24][0] = 8'h24;
frames[16][24][1] = 8'h6d;
frames[16][24][2] = 8'h6d;
frames[16][24][3] = 8'h6d;
frames[16][24][4] = 8'h48;
frames[16][24][5] = 8'h44;
frames[16][24][6] = 8'h6d;
frames[16][24][7] = 8'hb1;
frames[16][24][8] = 8'hd6;
frames[16][24][9] = 8'hda;
frames[16][24][10] = 8'hd6;
frames[16][24][11] = 8'hb1;
frames[16][24][12] = 8'hb1;
frames[16][24][13] = 8'h88;
frames[16][24][14] = 8'h8c;
frames[16][24][15] = 8'hb1;
frames[16][24][16] = 8'hb1;
frames[16][24][17] = 8'hd5;
frames[16][24][18] = 8'hd6;
frames[16][24][19] = 8'hd6;
frames[16][24][20] = 8'hb6;
frames[16][24][21] = 8'hb1;
frames[16][24][22] = 8'hb1;
frames[16][24][23] = 8'hb1;
frames[16][24][24] = 8'h6d;
frames[16][24][25] = 8'h44;
frames[16][24][26] = 8'h24;
frames[16][24][27] = 8'h24;
frames[16][24][28] = 8'h24;
frames[16][24][29] = 8'h24;
frames[16][24][30] = 8'h24;
frames[16][24][31] = 8'h48;
frames[16][24][32] = 8'h48;
frames[16][24][33] = 8'h48;
frames[16][24][34] = 8'h44;
frames[16][24][35] = 8'h69;
frames[16][24][36] = 8'hd6;
frames[16][24][37] = 8'hda;
frames[16][24][38] = 8'hd6;
frames[16][24][39] = 8'hb6;
frames[16][25][0] = 8'h44;
frames[16][25][1] = 8'h8d;
frames[16][25][2] = 8'h6d;
frames[16][25][3] = 8'h69;
frames[16][25][4] = 8'h48;
frames[16][25][5] = 8'h24;
frames[16][25][6] = 8'h20;
frames[16][25][7] = 8'h24;
frames[16][25][8] = 8'h49;
frames[16][25][9] = 8'h6d;
frames[16][25][10] = 8'h8d;
frames[16][25][11] = 8'h8d;
frames[16][25][12] = 8'h8d;
frames[16][25][13] = 8'h8d;
frames[16][25][14] = 8'h8d;
frames[16][25][15] = 8'h8d;
frames[16][25][16] = 8'h6d;
frames[16][25][17] = 8'h8d;
frames[16][25][18] = 8'h6d;
frames[16][25][19] = 8'h68;
frames[16][25][20] = 8'h48;
frames[16][25][21] = 8'h48;
frames[16][25][22] = 8'h48;
frames[16][25][23] = 8'h44;
frames[16][25][24] = 8'h44;
frames[16][25][25] = 8'h44;
frames[16][25][26] = 8'h48;
frames[16][25][27] = 8'h48;
frames[16][25][28] = 8'h49;
frames[16][25][29] = 8'h49;
frames[16][25][30] = 8'h49;
frames[16][25][31] = 8'h48;
frames[16][25][32] = 8'h48;
frames[16][25][33] = 8'h44;
frames[16][25][34] = 8'h44;
frames[16][25][35] = 8'hb2;
frames[16][25][36] = 8'hda;
frames[16][25][37] = 8'hd6;
frames[16][25][38] = 8'hd6;
frames[16][25][39] = 8'hb6;
frames[16][26][0] = 8'h48;
frames[16][26][1] = 8'h6d;
frames[16][26][2] = 8'h69;
frames[16][26][3] = 8'h48;
frames[16][26][4] = 8'h48;
frames[16][26][5] = 8'h44;
frames[16][26][6] = 8'h24;
frames[16][26][7] = 8'h24;
frames[16][26][8] = 8'h24;
frames[16][26][9] = 8'h24;
frames[16][26][10] = 8'h24;
frames[16][26][11] = 8'h44;
frames[16][26][12] = 8'h44;
frames[16][26][13] = 8'h44;
frames[16][26][14] = 8'h44;
frames[16][26][15] = 8'h44;
frames[16][26][16] = 8'h44;
frames[16][26][17] = 8'h24;
frames[16][26][18] = 8'h44;
frames[16][26][19] = 8'h44;
frames[16][26][20] = 8'h44;
frames[16][26][21] = 8'h44;
frames[16][26][22] = 8'h44;
frames[16][26][23] = 8'h48;
frames[16][26][24] = 8'h49;
frames[16][26][25] = 8'h48;
frames[16][26][26] = 8'h44;
frames[16][26][27] = 8'h44;
frames[16][26][28] = 8'h44;
frames[16][26][29] = 8'h44;
frames[16][26][30] = 8'h44;
frames[16][26][31] = 8'h44;
frames[16][26][32] = 8'h24;
frames[16][26][33] = 8'h24;
frames[16][26][34] = 8'h44;
frames[16][26][35] = 8'h8d;
frames[16][26][36] = 8'hd6;
frames[16][26][37] = 8'hb6;
frames[16][26][38] = 8'hb6;
frames[16][26][39] = 8'hb2;
frames[16][27][0] = 8'h24;
frames[16][27][1] = 8'h24;
frames[16][27][2] = 8'h44;
frames[16][27][3] = 8'h24;
frames[16][27][4] = 8'h44;
frames[16][27][5] = 8'h24;
frames[16][27][6] = 8'h44;
frames[16][27][7] = 8'h44;
frames[16][27][8] = 8'h44;
frames[16][27][9] = 8'h24;
frames[16][27][10] = 8'h24;
frames[16][27][11] = 8'h24;
frames[16][27][12] = 8'h24;
frames[16][27][13] = 8'h24;
frames[16][27][14] = 8'h24;
frames[16][27][15] = 8'h24;
frames[16][27][16] = 8'h24;
frames[16][27][17] = 8'h24;
frames[16][27][18] = 8'h24;
frames[16][27][19] = 8'h24;
frames[16][27][20] = 8'h24;
frames[16][27][21] = 8'h24;
frames[16][27][22] = 8'h24;
frames[16][27][23] = 8'h24;
frames[16][27][24] = 8'h24;
frames[16][27][25] = 8'h24;
frames[16][27][26] = 8'h24;
frames[16][27][27] = 8'h24;
frames[16][27][28] = 8'h24;
frames[16][27][29] = 8'h24;
frames[16][27][30] = 8'h24;
frames[16][27][31] = 8'h24;
frames[16][27][32] = 8'h24;
frames[16][27][33] = 8'h44;
frames[16][27][34] = 8'h44;
frames[16][27][35] = 8'h68;
frames[16][27][36] = 8'hb6;
frames[16][27][37] = 8'hb2;
frames[16][27][38] = 8'hb2;
frames[16][27][39] = 8'hb1;
frames[16][28][0] = 8'h24;
frames[16][28][1] = 8'h24;
frames[16][28][2] = 8'h24;
frames[16][28][3] = 8'h24;
frames[16][28][4] = 8'h44;
frames[16][28][5] = 8'h24;
frames[16][28][6] = 8'h44;
frames[16][28][7] = 8'h44;
frames[16][28][8] = 8'h44;
frames[16][28][9] = 8'h44;
frames[16][28][10] = 8'h44;
frames[16][28][11] = 8'h24;
frames[16][28][12] = 8'h24;
frames[16][28][13] = 8'h24;
frames[16][28][14] = 8'h44;
frames[16][28][15] = 8'h44;
frames[16][28][16] = 8'h44;
frames[16][28][17] = 8'h44;
frames[16][28][18] = 8'h44;
frames[16][28][19] = 8'h44;
frames[16][28][20] = 8'h44;
frames[16][28][21] = 8'h44;
frames[16][28][22] = 8'h44;
frames[16][28][23] = 8'h44;
frames[16][28][24] = 8'h44;
frames[16][28][25] = 8'h44;
frames[16][28][26] = 8'h44;
frames[16][28][27] = 8'h44;
frames[16][28][28] = 8'h44;
frames[16][28][29] = 8'h44;
frames[16][28][30] = 8'h44;
frames[16][28][31] = 8'h44;
frames[16][28][32] = 8'h44;
frames[16][28][33] = 8'h44;
frames[16][28][34] = 8'h44;
frames[16][28][35] = 8'h68;
frames[16][28][36] = 8'hb2;
frames[16][28][37] = 8'hb2;
frames[16][28][38] = 8'hb1;
frames[16][28][39] = 8'hb1;
frames[16][29][0] = 8'h44;
frames[16][29][1] = 8'h44;
frames[16][29][2] = 8'h44;
frames[16][29][3] = 8'h44;
frames[16][29][4] = 8'h44;
frames[16][29][5] = 8'h44;
frames[16][29][6] = 8'h44;
frames[16][29][7] = 8'h44;
frames[16][29][8] = 8'h44;
frames[16][29][9] = 8'h44;
frames[16][29][10] = 8'h44;
frames[16][29][11] = 8'h44;
frames[16][29][12] = 8'h44;
frames[16][29][13] = 8'h44;
frames[16][29][14] = 8'h44;
frames[16][29][15] = 8'h44;
frames[16][29][16] = 8'h44;
frames[16][29][17] = 8'h64;
frames[16][29][18] = 8'h64;
frames[16][29][19] = 8'h44;
frames[16][29][20] = 8'h64;
frames[16][29][21] = 8'h64;
frames[16][29][22] = 8'h64;
frames[16][29][23] = 8'h64;
frames[16][29][24] = 8'h64;
frames[16][29][25] = 8'h64;
frames[16][29][26] = 8'h64;
frames[16][29][27] = 8'h64;
frames[16][29][28] = 8'h64;
frames[16][29][29] = 8'h64;
frames[16][29][30] = 8'h64;
frames[16][29][31] = 8'h64;
frames[16][29][32] = 8'h68;
frames[16][29][33] = 8'h68;
frames[16][29][34] = 8'h68;
frames[16][29][35] = 8'h68;
frames[16][29][36] = 8'h91;
frames[16][29][37] = 8'hb1;
frames[16][29][38] = 8'h8d;
frames[16][29][39] = 8'h8d;
frames[17][0][0] = 8'hff;
frames[17][0][1] = 8'hfa;
frames[17][0][2] = 8'hb1;
frames[17][0][3] = 8'h48;
frames[17][0][4] = 8'h64;
frames[17][0][5] = 8'h68;
frames[17][0][6] = 8'h69;
frames[17][0][7] = 8'h48;
frames[17][0][8] = 8'h44;
frames[17][0][9] = 8'h48;
frames[17][0][10] = 8'h48;
frames[17][0][11] = 8'h6d;
frames[17][0][12] = 8'h69;
frames[17][0][13] = 8'h48;
frames[17][0][14] = 8'h44;
frames[17][0][15] = 8'h44;
frames[17][0][16] = 8'h44;
frames[17][0][17] = 8'h44;
frames[17][0][18] = 8'h24;
frames[17][0][19] = 8'h48;
frames[17][0][20] = 8'h48;
frames[17][0][21] = 8'h48;
frames[17][0][22] = 8'h44;
frames[17][0][23] = 8'h48;
frames[17][0][24] = 8'h49;
frames[17][0][25] = 8'h44;
frames[17][0][26] = 8'h44;
frames[17][0][27] = 8'h49;
frames[17][0][28] = 8'h49;
frames[17][0][29] = 8'h48;
frames[17][0][30] = 8'h24;
frames[17][0][31] = 8'h44;
frames[17][0][32] = 8'h44;
frames[17][0][33] = 8'h24;
frames[17][0][34] = 8'h44;
frames[17][0][35] = 8'h24;
frames[17][0][36] = 8'h00;
frames[17][0][37] = 8'h48;
frames[17][0][38] = 8'h24;
frames[17][0][39] = 8'h00;
frames[17][1][0] = 8'h8d;
frames[17][1][1] = 8'h88;
frames[17][1][2] = 8'h69;
frames[17][1][3] = 8'h8d;
frames[17][1][4] = 8'h68;
frames[17][1][5] = 8'h68;
frames[17][1][6] = 8'h68;
frames[17][1][7] = 8'h48;
frames[17][1][8] = 8'h44;
frames[17][1][9] = 8'h44;
frames[17][1][10] = 8'h48;
frames[17][1][11] = 8'h44;
frames[17][1][12] = 8'h44;
frames[17][1][13] = 8'h44;
frames[17][1][14] = 8'h44;
frames[17][1][15] = 8'h44;
frames[17][1][16] = 8'h44;
frames[17][1][17] = 8'h44;
frames[17][1][18] = 8'h44;
frames[17][1][19] = 8'h48;
frames[17][1][20] = 8'h48;
frames[17][1][21] = 8'h44;
frames[17][1][22] = 8'h44;
frames[17][1][23] = 8'h69;
frames[17][1][24] = 8'h48;
frames[17][1][25] = 8'h44;
frames[17][1][26] = 8'h44;
frames[17][1][27] = 8'h49;
frames[17][1][28] = 8'h69;
frames[17][1][29] = 8'h48;
frames[17][1][30] = 8'h44;
frames[17][1][31] = 8'h48;
frames[17][1][32] = 8'h48;
frames[17][1][33] = 8'h48;
frames[17][1][34] = 8'h48;
frames[17][1][35] = 8'h24;
frames[17][1][36] = 8'h49;
frames[17][1][37] = 8'hb6;
frames[17][1][38] = 8'hb6;
frames[17][1][39] = 8'h24;
frames[17][2][0] = 8'h68;
frames[17][2][1] = 8'h8d;
frames[17][2][2] = 8'h8d;
frames[17][2][3] = 8'h8d;
frames[17][2][4] = 8'h68;
frames[17][2][5] = 8'h48;
frames[17][2][6] = 8'h44;
frames[17][2][7] = 8'h48;
frames[17][2][8] = 8'h44;
frames[17][2][9] = 8'h48;
frames[17][2][10] = 8'h48;
frames[17][2][11] = 8'h44;
frames[17][2][12] = 8'h44;
frames[17][2][13] = 8'h48;
frames[17][2][14] = 8'h44;
frames[17][2][15] = 8'h44;
frames[17][2][16] = 8'h44;
frames[17][2][17] = 8'h44;
frames[17][2][18] = 8'h24;
frames[17][2][19] = 8'h44;
frames[17][2][20] = 8'h48;
frames[17][2][21] = 8'h44;
frames[17][2][22] = 8'h48;
frames[17][2][23] = 8'h69;
frames[17][2][24] = 8'h49;
frames[17][2][25] = 8'h48;
frames[17][2][26] = 8'h48;
frames[17][2][27] = 8'h69;
frames[17][2][28] = 8'h48;
frames[17][2][29] = 8'h48;
frames[17][2][30] = 8'h44;
frames[17][2][31] = 8'h44;
frames[17][2][32] = 8'h24;
frames[17][2][33] = 8'h24;
frames[17][2][34] = 8'h24;
frames[17][2][35] = 8'h24;
frames[17][2][36] = 8'h92;
frames[17][2][37] = 8'h6d;
frames[17][2][38] = 8'h4d;
frames[17][2][39] = 8'h6e;
frames[17][3][0] = 8'h69;
frames[17][3][1] = 8'h69;
frames[17][3][2] = 8'h44;
frames[17][3][3] = 8'h44;
frames[17][3][4] = 8'h44;
frames[17][3][5] = 8'h24;
frames[17][3][6] = 8'h44;
frames[17][3][7] = 8'h44;
frames[17][3][8] = 8'h44;
frames[17][3][9] = 8'h48;
frames[17][3][10] = 8'h48;
frames[17][3][11] = 8'h44;
frames[17][3][12] = 8'h44;
frames[17][3][13] = 8'h44;
frames[17][3][14] = 8'h44;
frames[17][3][15] = 8'h44;
frames[17][3][16] = 8'h48;
frames[17][3][17] = 8'h44;
frames[17][3][18] = 8'h48;
frames[17][3][19] = 8'h48;
frames[17][3][20] = 8'h48;
frames[17][3][21] = 8'h48;
frames[17][3][22] = 8'h48;
frames[17][3][23] = 8'h49;
frames[17][3][24] = 8'h48;
frames[17][3][25] = 8'h48;
frames[17][3][26] = 8'h44;
frames[17][3][27] = 8'h24;
frames[17][3][28] = 8'h24;
frames[17][3][29] = 8'h44;
frames[17][3][30] = 8'h24;
frames[17][3][31] = 8'h24;
frames[17][3][32] = 8'h24;
frames[17][3][33] = 8'h24;
frames[17][3][34] = 8'h24;
frames[17][3][35] = 8'h48;
frames[17][3][36] = 8'h92;
frames[17][3][37] = 8'h6d;
frames[17][3][38] = 8'h49;
frames[17][3][39] = 8'h72;
frames[17][4][0] = 8'h48;
frames[17][4][1] = 8'h68;
frames[17][4][2] = 8'h44;
frames[17][4][3] = 8'h44;
frames[17][4][4] = 8'h44;
frames[17][4][5] = 8'h48;
frames[17][4][6] = 8'h68;
frames[17][4][7] = 8'h69;
frames[17][4][8] = 8'h69;
frames[17][4][9] = 8'h69;
frames[17][4][10] = 8'h68;
frames[17][4][11] = 8'h48;
frames[17][4][12] = 8'h48;
frames[17][4][13] = 8'h49;
frames[17][4][14] = 8'h49;
frames[17][4][15] = 8'h49;
frames[17][4][16] = 8'h49;
frames[17][4][17] = 8'h48;
frames[17][4][18] = 8'h49;
frames[17][4][19] = 8'h48;
frames[17][4][20] = 8'h44;
frames[17][4][21] = 8'h48;
frames[17][4][22] = 8'h44;
frames[17][4][23] = 8'h44;
frames[17][4][24] = 8'h44;
frames[17][4][25] = 8'h44;
frames[17][4][26] = 8'h24;
frames[17][4][27] = 8'h24;
frames[17][4][28] = 8'h24;
frames[17][4][29] = 8'h24;
frames[17][4][30] = 8'h24;
frames[17][4][31] = 8'h24;
frames[17][4][32] = 8'h24;
frames[17][4][33] = 8'h24;
frames[17][4][34] = 8'h24;
frames[17][4][35] = 8'h24;
frames[17][4][36] = 8'h92;
frames[17][4][37] = 8'h6d;
frames[17][4][38] = 8'h6e;
frames[17][4][39] = 8'h6e;
frames[17][5][0] = 8'h48;
frames[17][5][1] = 8'h69;
frames[17][5][2] = 8'h69;
frames[17][5][3] = 8'h69;
frames[17][5][4] = 8'h6d;
frames[17][5][5] = 8'h6d;
frames[17][5][6] = 8'h6d;
frames[17][5][7] = 8'h6d;
frames[17][5][8] = 8'h8d;
frames[17][5][9] = 8'h8d;
frames[17][5][10] = 8'h6d;
frames[17][5][11] = 8'h48;
frames[17][5][12] = 8'h48;
frames[17][5][13] = 8'h48;
frames[17][5][14] = 8'h48;
frames[17][5][15] = 8'h48;
frames[17][5][16] = 8'h48;
frames[17][5][17] = 8'h28;
frames[17][5][18] = 8'h44;
frames[17][5][19] = 8'h44;
frames[17][5][20] = 8'h44;
frames[17][5][21] = 8'h44;
frames[17][5][22] = 8'h44;
frames[17][5][23] = 8'h44;
frames[17][5][24] = 8'h24;
frames[17][5][25] = 8'h24;
frames[17][5][26] = 8'h24;
frames[17][5][27] = 8'h24;
frames[17][5][28] = 8'h24;
frames[17][5][29] = 8'h24;
frames[17][5][30] = 8'h24;
frames[17][5][31] = 8'h24;
frames[17][5][32] = 8'h24;
frames[17][5][33] = 8'h24;
frames[17][5][34] = 8'h24;
frames[17][5][35] = 8'h24;
frames[17][5][36] = 8'h49;
frames[17][5][37] = 8'h92;
frames[17][5][38] = 8'h92;
frames[17][5][39] = 8'h24;
frames[17][6][0] = 8'h6d;
frames[17][6][1] = 8'h6d;
frames[17][6][2] = 8'h6d;
frames[17][6][3] = 8'h6d;
frames[17][6][4] = 8'h6d;
frames[17][6][5] = 8'h6d;
frames[17][6][6] = 8'h69;
frames[17][6][7] = 8'h69;
frames[17][6][8] = 8'h6d;
frames[17][6][9] = 8'h6d;
frames[17][6][10] = 8'h69;
frames[17][6][11] = 8'h24;
frames[17][6][12] = 8'h24;
frames[17][6][13] = 8'h24;
frames[17][6][14] = 8'h24;
frames[17][6][15] = 8'h28;
frames[17][6][16] = 8'h28;
frames[17][6][17] = 8'h48;
frames[17][6][18] = 8'h48;
frames[17][6][19] = 8'h44;
frames[17][6][20] = 8'h44;
frames[17][6][21] = 8'h44;
frames[17][6][22] = 8'h44;
frames[17][6][23] = 8'h44;
frames[17][6][24] = 8'h24;
frames[17][6][25] = 8'h24;
frames[17][6][26] = 8'h24;
frames[17][6][27] = 8'h24;
frames[17][6][28] = 8'h24;
frames[17][6][29] = 8'h24;
frames[17][6][30] = 8'h24;
frames[17][6][31] = 8'h24;
frames[17][6][32] = 8'h24;
frames[17][6][33] = 8'h24;
frames[17][6][34] = 8'h24;
frames[17][6][35] = 8'h24;
frames[17][6][36] = 8'h24;
frames[17][6][37] = 8'h24;
frames[17][6][38] = 8'h24;
frames[17][6][39] = 8'h24;
frames[17][7][0] = 8'h49;
frames[17][7][1] = 8'h6d;
frames[17][7][2] = 8'h6d;
frames[17][7][3] = 8'h6d;
frames[17][7][4] = 8'h6d;
frames[17][7][5] = 8'h6d;
frames[17][7][6] = 8'h6d;
frames[17][7][7] = 8'h6d;
frames[17][7][8] = 8'h6d;
frames[17][7][9] = 8'h6d;
frames[17][7][10] = 8'h48;
frames[17][7][11] = 8'h24;
frames[17][7][12] = 8'h24;
frames[17][7][13] = 8'h24;
frames[17][7][14] = 8'h24;
frames[17][7][15] = 8'h44;
frames[17][7][16] = 8'h48;
frames[17][7][17] = 8'h48;
frames[17][7][18] = 8'h44;
frames[17][7][19] = 8'h44;
frames[17][7][20] = 8'h44;
frames[17][7][21] = 8'h44;
frames[17][7][22] = 8'h44;
frames[17][7][23] = 8'h44;
frames[17][7][24] = 8'h24;
frames[17][7][25] = 8'h24;
frames[17][7][26] = 8'h24;
frames[17][7][27] = 8'h24;
frames[17][7][28] = 8'h24;
frames[17][7][29] = 8'h24;
frames[17][7][30] = 8'h24;
frames[17][7][31] = 8'h24;
frames[17][7][32] = 8'h24;
frames[17][7][33] = 8'h24;
frames[17][7][34] = 8'h24;
frames[17][7][35] = 8'h24;
frames[17][7][36] = 8'h24;
frames[17][7][37] = 8'h24;
frames[17][7][38] = 8'h24;
frames[17][7][39] = 8'h24;
frames[17][8][0] = 8'h24;
frames[17][8][1] = 8'h24;
frames[17][8][2] = 8'h24;
frames[17][8][3] = 8'h48;
frames[17][8][4] = 8'h48;
frames[17][8][5] = 8'h49;
frames[17][8][6] = 8'h49;
frames[17][8][7] = 8'h6d;
frames[17][8][8] = 8'h6d;
frames[17][8][9] = 8'h6d;
frames[17][8][10] = 8'h44;
frames[17][8][11] = 8'h24;
frames[17][8][12] = 8'h24;
frames[17][8][13] = 8'h44;
frames[17][8][14] = 8'h24;
frames[17][8][15] = 8'h44;
frames[17][8][16] = 8'h24;
frames[17][8][17] = 8'h24;
frames[17][8][18] = 8'h44;
frames[17][8][19] = 8'h44;
frames[17][8][20] = 8'h44;
frames[17][8][21] = 8'h44;
frames[17][8][22] = 8'h44;
frames[17][8][23] = 8'h44;
frames[17][8][24] = 8'h24;
frames[17][8][25] = 8'h24;
frames[17][8][26] = 8'h24;
frames[17][8][27] = 8'h24;
frames[17][8][28] = 8'h24;
frames[17][8][29] = 8'h24;
frames[17][8][30] = 8'h24;
frames[17][8][31] = 8'h24;
frames[17][8][32] = 8'h24;
frames[17][8][33] = 8'h24;
frames[17][8][34] = 8'h24;
frames[17][8][35] = 8'h24;
frames[17][8][36] = 8'h24;
frames[17][8][37] = 8'h24;
frames[17][8][38] = 8'h24;
frames[17][8][39] = 8'h24;
frames[17][9][0] = 8'h24;
frames[17][9][1] = 8'h24;
frames[17][9][2] = 8'h24;
frames[17][9][3] = 8'h48;
frames[17][9][4] = 8'h6d;
frames[17][9][5] = 8'h92;
frames[17][9][6] = 8'hb6;
frames[17][9][7] = 8'hda;
frames[17][9][8] = 8'hdb;
frames[17][9][9] = 8'hb6;
frames[17][9][10] = 8'h24;
frames[17][9][11] = 8'h24;
frames[17][9][12] = 8'h24;
frames[17][9][13] = 8'h24;
frames[17][9][14] = 8'h24;
frames[17][9][15] = 8'h44;
frames[17][9][16] = 8'h24;
frames[17][9][17] = 8'h44;
frames[17][9][18] = 8'h44;
frames[17][9][19] = 8'h44;
frames[17][9][20] = 8'h44;
frames[17][9][21] = 8'h44;
frames[17][9][22] = 8'h44;
frames[17][9][23] = 8'h44;
frames[17][9][24] = 8'h44;
frames[17][9][25] = 8'h44;
frames[17][9][26] = 8'h24;
frames[17][9][27] = 8'h24;
frames[17][9][28] = 8'h24;
frames[17][9][29] = 8'h24;
frames[17][9][30] = 8'h24;
frames[17][9][31] = 8'h48;
frames[17][9][32] = 8'h48;
frames[17][9][33] = 8'h24;
frames[17][9][34] = 8'h24;
frames[17][9][35] = 8'h24;
frames[17][9][36] = 8'h24;
frames[17][9][37] = 8'h24;
frames[17][9][38] = 8'h24;
frames[17][9][39] = 8'h24;
frames[17][10][0] = 8'h92;
frames[17][10][1] = 8'hb6;
frames[17][10][2] = 8'hb6;
frames[17][10][3] = 8'hdb;
frames[17][10][4] = 8'hdb;
frames[17][10][5] = 8'hda;
frames[17][10][6] = 8'hda;
frames[17][10][7] = 8'hb6;
frames[17][10][8] = 8'hda;
frames[17][10][9] = 8'h6d;
frames[17][10][10] = 8'h24;
frames[17][10][11] = 8'h24;
frames[17][10][12] = 8'h24;
frames[17][10][13] = 8'h24;
frames[17][10][14] = 8'h24;
frames[17][10][15] = 8'h24;
frames[17][10][16] = 8'h24;
frames[17][10][17] = 8'h44;
frames[17][10][18] = 8'h44;
frames[17][10][19] = 8'h44;
frames[17][10][20] = 8'h44;
frames[17][10][21] = 8'h44;
frames[17][10][22] = 8'h44;
frames[17][10][23] = 8'h44;
frames[17][10][24] = 8'h24;
frames[17][10][25] = 8'h24;
frames[17][10][26] = 8'h24;
frames[17][10][27] = 8'h48;
frames[17][10][28] = 8'h91;
frames[17][10][29] = 8'hda;
frames[17][10][30] = 8'hdb;
frames[17][10][31] = 8'hff;
frames[17][10][32] = 8'hff;
frames[17][10][33] = 8'hdb;
frames[17][10][34] = 8'h92;
frames[17][10][35] = 8'h48;
frames[17][10][36] = 8'h24;
frames[17][10][37] = 8'h24;
frames[17][10][38] = 8'h24;
frames[17][10][39] = 8'h24;
frames[17][11][0] = 8'hb6;
frames[17][11][1] = 8'hb6;
frames[17][11][2] = 8'hb6;
frames[17][11][3] = 8'hb6;
frames[17][11][4] = 8'hb6;
frames[17][11][5] = 8'hb6;
frames[17][11][6] = 8'hda;
frames[17][11][7] = 8'hdb;
frames[17][11][8] = 8'hdb;
frames[17][11][9] = 8'h48;
frames[17][11][10] = 8'h24;
frames[17][11][11] = 8'h24;
frames[17][11][12] = 8'h24;
frames[17][11][13] = 8'h24;
frames[17][11][14] = 8'h24;
frames[17][11][15] = 8'h44;
frames[17][11][16] = 8'h44;
frames[17][11][17] = 8'h44;
frames[17][11][18] = 8'h24;
frames[17][11][19] = 8'h24;
frames[17][11][20] = 8'h44;
frames[17][11][21] = 8'h44;
frames[17][11][22] = 8'h24;
frames[17][11][23] = 8'h44;
frames[17][11][24] = 8'h69;
frames[17][11][25] = 8'h91;
frames[17][11][26] = 8'hb6;
frames[17][11][27] = 8'hfb;
frames[17][11][28] = 8'hff;
frames[17][11][29] = 8'hff;
frames[17][11][30] = 8'hff;
frames[17][11][31] = 8'hff;
frames[17][11][32] = 8'hff;
frames[17][11][33] = 8'hff;
frames[17][11][34] = 8'hff;
frames[17][11][35] = 8'hff;
frames[17][11][36] = 8'h92;
frames[17][11][37] = 8'h24;
frames[17][11][38] = 8'h24;
frames[17][11][39] = 8'h24;
frames[17][12][0] = 8'hb6;
frames[17][12][1] = 8'hb6;
frames[17][12][2] = 8'hda;
frames[17][12][3] = 8'hdb;
frames[17][12][4] = 8'hdf;
frames[17][12][5] = 8'hdf;
frames[17][12][6] = 8'hff;
frames[17][12][7] = 8'hff;
frames[17][12][8] = 8'hb6;
frames[17][12][9] = 8'h24;
frames[17][12][10] = 8'h24;
frames[17][12][11] = 8'h24;
frames[17][12][12] = 8'h24;
frames[17][12][13] = 8'h24;
frames[17][12][14] = 8'h24;
frames[17][12][15] = 8'h24;
frames[17][12][16] = 8'h44;
frames[17][12][17] = 8'h44;
frames[17][12][18] = 8'h24;
frames[17][12][19] = 8'h24;
frames[17][12][20] = 8'h24;
frames[17][12][21] = 8'h24;
frames[17][12][22] = 8'h92;
frames[17][12][23] = 8'hfb;
frames[17][12][24] = 8'hff;
frames[17][12][25] = 8'hff;
frames[17][12][26] = 8'hff;
frames[17][12][27] = 8'hff;
frames[17][12][28] = 8'hff;
frames[17][12][29] = 8'hff;
frames[17][12][30] = 8'hff;
frames[17][12][31] = 8'hff;
frames[17][12][32] = 8'hff;
frames[17][12][33] = 8'hff;
frames[17][12][34] = 8'hff;
frames[17][12][35] = 8'hff;
frames[17][12][36] = 8'hff;
frames[17][12][37] = 8'hdb;
frames[17][12][38] = 8'h48;
frames[17][12][39] = 8'h00;
frames[17][13][0] = 8'hdb;
frames[17][13][1] = 8'hdb;
frames[17][13][2] = 8'hdf;
frames[17][13][3] = 8'hdf;
frames[17][13][4] = 8'hff;
frames[17][13][5] = 8'hff;
frames[17][13][6] = 8'hff;
frames[17][13][7] = 8'hff;
frames[17][13][8] = 8'h91;
frames[17][13][9] = 8'h24;
frames[17][13][10] = 8'h24;
frames[17][13][11] = 8'h24;
frames[17][13][12] = 8'h24;
frames[17][13][13] = 8'h24;
frames[17][13][14] = 8'h24;
frames[17][13][15] = 8'h24;
frames[17][13][16] = 8'h24;
frames[17][13][17] = 8'h24;
frames[17][13][18] = 8'h24;
frames[17][13][19] = 8'h24;
frames[17][13][20] = 8'h24;
frames[17][13][21] = 8'h6d;
frames[17][13][22] = 8'hff;
frames[17][13][23] = 8'hff;
frames[17][13][24] = 8'hff;
frames[17][13][25] = 8'hff;
frames[17][13][26] = 8'hff;
frames[17][13][27] = 8'hff;
frames[17][13][28] = 8'hff;
frames[17][13][29] = 8'hff;
frames[17][13][30] = 8'hff;
frames[17][13][31] = 8'hff;
frames[17][13][32] = 8'hff;
frames[17][13][33] = 8'hff;
frames[17][13][34] = 8'hff;
frames[17][13][35] = 8'hff;
frames[17][13][36] = 8'hff;
frames[17][13][37] = 8'hff;
frames[17][13][38] = 8'hda;
frames[17][13][39] = 8'h24;
frames[17][14][0] = 8'hdb;
frames[17][14][1] = 8'hdb;
frames[17][14][2] = 8'hdf;
frames[17][14][3] = 8'hdf;
frames[17][14][4] = 8'hdb;
frames[17][14][5] = 8'hdb;
frames[17][14][6] = 8'hb6;
frames[17][14][7] = 8'h96;
frames[17][14][8] = 8'h48;
frames[17][14][9] = 8'h24;
frames[17][14][10] = 8'h24;
frames[17][14][11] = 8'h24;
frames[17][14][12] = 8'h24;
frames[17][14][13] = 8'h24;
frames[17][14][14] = 8'h24;
frames[17][14][15] = 8'h24;
frames[17][14][16] = 8'h24;
frames[17][14][17] = 8'h24;
frames[17][14][18] = 8'h24;
frames[17][14][19] = 8'h24;
frames[17][14][20] = 8'h24;
frames[17][14][21] = 8'hb6;
frames[17][14][22] = 8'hff;
frames[17][14][23] = 8'hff;
frames[17][14][24] = 8'hff;
frames[17][14][25] = 8'hff;
frames[17][14][26] = 8'hff;
frames[17][14][27] = 8'hff;
frames[17][14][28] = 8'hff;
frames[17][14][29] = 8'hff;
frames[17][14][30] = 8'hff;
frames[17][14][31] = 8'hff;
frames[17][14][32] = 8'hff;
frames[17][14][33] = 8'hff;
frames[17][14][34] = 8'hff;
frames[17][14][35] = 8'hff;
frames[17][14][36] = 8'hff;
frames[17][14][37] = 8'hff;
frames[17][14][38] = 8'hff;
frames[17][14][39] = 8'h49;
frames[17][15][0] = 8'hba;
frames[17][15][1] = 8'hb6;
frames[17][15][2] = 8'h91;
frames[17][15][3] = 8'h6d;
frames[17][15][4] = 8'h49;
frames[17][15][5] = 8'h24;
frames[17][15][6] = 8'h24;
frames[17][15][7] = 8'h24;
frames[17][15][8] = 8'h24;
frames[17][15][9] = 8'h24;
frames[17][15][10] = 8'h24;
frames[17][15][11] = 8'h24;
frames[17][15][12] = 8'h24;
frames[17][15][13] = 8'h24;
frames[17][15][14] = 8'h24;
frames[17][15][15] = 8'h24;
frames[17][15][16] = 8'h24;
frames[17][15][17] = 8'h24;
frames[17][15][18] = 8'h24;
frames[17][15][19] = 8'h24;
frames[17][15][20] = 8'h24;
frames[17][15][21] = 8'h24;
frames[17][15][22] = 8'hd6;
frames[17][15][23] = 8'hff;
frames[17][15][24] = 8'hff;
frames[17][15][25] = 8'hff;
frames[17][15][26] = 8'hff;
frames[17][15][27] = 8'hff;
frames[17][15][28] = 8'hff;
frames[17][15][29] = 8'hff;
frames[17][15][30] = 8'hff;
frames[17][15][31] = 8'hff;
frames[17][15][32] = 8'hff;
frames[17][15][33] = 8'hff;
frames[17][15][34] = 8'hff;
frames[17][15][35] = 8'hff;
frames[17][15][36] = 8'hff;
frames[17][15][37] = 8'hff;
frames[17][15][38] = 8'hb6;
frames[17][15][39] = 8'h24;
frames[17][16][0] = 8'h44;
frames[17][16][1] = 8'h24;
frames[17][16][2] = 8'h24;
frames[17][16][3] = 8'h24;
frames[17][16][4] = 8'h24;
frames[17][16][5] = 8'h24;
frames[17][16][6] = 8'h24;
frames[17][16][7] = 8'h24;
frames[17][16][8] = 8'h24;
frames[17][16][9] = 8'h24;
frames[17][16][10] = 8'h24;
frames[17][16][11] = 8'h24;
frames[17][16][12] = 8'h24;
frames[17][16][13] = 8'h24;
frames[17][16][14] = 8'h24;
frames[17][16][15] = 8'h24;
frames[17][16][16] = 8'h24;
frames[17][16][17] = 8'h24;
frames[17][16][18] = 8'h24;
frames[17][16][19] = 8'h24;
frames[17][16][20] = 8'h24;
frames[17][16][21] = 8'h00;
frames[17][16][22] = 8'h64;
frames[17][16][23] = 8'h8d;
frames[17][16][24] = 8'hb2;
frames[17][16][25] = 8'hd6;
frames[17][16][26] = 8'hfb;
frames[17][16][27] = 8'hff;
frames[17][16][28] = 8'hff;
frames[17][16][29] = 8'hff;
frames[17][16][30] = 8'hff;
frames[17][16][31] = 8'hff;
frames[17][16][32] = 8'hff;
frames[17][16][33] = 8'hff;
frames[17][16][34] = 8'hfa;
frames[17][16][35] = 8'hd6;
frames[17][16][36] = 8'hb1;
frames[17][16][37] = 8'h8d;
frames[17][16][38] = 8'h49;
frames[17][16][39] = 8'h00;
frames[17][17][0] = 8'h49;
frames[17][17][1] = 8'h44;
frames[17][17][2] = 8'h24;
frames[17][17][3] = 8'h24;
frames[17][17][4] = 8'h24;
frames[17][17][5] = 8'h24;
frames[17][17][6] = 8'h24;
frames[17][17][7] = 8'h24;
frames[17][17][8] = 8'h24;
frames[17][17][9] = 8'h24;
frames[17][17][10] = 8'h24;
frames[17][17][11] = 8'h24;
frames[17][17][12] = 8'h24;
frames[17][17][13] = 8'h24;
frames[17][17][14] = 8'h24;
frames[17][17][15] = 8'h24;
frames[17][17][16] = 8'h24;
frames[17][17][17] = 8'h24;
frames[17][17][18] = 8'h24;
frames[17][17][19] = 8'h44;
frames[17][17][20] = 8'h44;
frames[17][17][21] = 8'h24;
frames[17][17][22] = 8'h20;
frames[17][17][23] = 8'h64;
frames[17][17][24] = 8'h89;
frames[17][17][25] = 8'h89;
frames[17][17][26] = 8'h88;
frames[17][17][27] = 8'had;
frames[17][17][28] = 8'hb1;
frames[17][17][29] = 8'hd6;
frames[17][17][30] = 8'hb1;
frames[17][17][31] = 8'hb1;
frames[17][17][32] = 8'hb1;
frames[17][17][33] = 8'h91;
frames[17][17][34] = 8'hb1;
frames[17][17][35] = 8'h8d;
frames[17][17][36] = 8'h64;
frames[17][17][37] = 8'h68;
frames[17][17][38] = 8'h24;
frames[17][17][39] = 8'h00;
frames[17][18][0] = 8'h24;
frames[17][18][1] = 8'h44;
frames[17][18][2] = 8'h49;
frames[17][18][3] = 8'h49;
frames[17][18][4] = 8'h44;
frames[17][18][5] = 8'h24;
frames[17][18][6] = 8'h24;
frames[17][18][7] = 8'h24;
frames[17][18][8] = 8'h24;
frames[17][18][9] = 8'h24;
frames[17][18][10] = 8'h24;
frames[17][18][11] = 8'h24;
frames[17][18][12] = 8'h24;
frames[17][18][13] = 8'h24;
frames[17][18][14] = 8'h24;
frames[17][18][15] = 8'h24;
frames[17][18][16] = 8'h24;
frames[17][18][17] = 8'h24;
frames[17][18][18] = 8'h44;
frames[17][18][19] = 8'h44;
frames[17][18][20] = 8'h24;
frames[17][18][21] = 8'h24;
frames[17][18][22] = 8'h24;
frames[17][18][23] = 8'h44;
frames[17][18][24] = 8'h44;
frames[17][18][25] = 8'h44;
frames[17][18][26] = 8'h44;
frames[17][18][27] = 8'h69;
frames[17][18][28] = 8'h8d;
frames[17][18][29] = 8'h8d;
frames[17][18][30] = 8'h8d;
frames[17][18][31] = 8'h8d;
frames[17][18][32] = 8'h91;
frames[17][18][33] = 8'h91;
frames[17][18][34] = 8'h8d;
frames[17][18][35] = 8'h69;
frames[17][18][36] = 8'h24;
frames[17][18][37] = 8'h20;
frames[17][18][38] = 8'h00;
frames[17][18][39] = 8'h04;
frames[17][19][0] = 8'h24;
frames[17][19][1] = 8'h24;
frames[17][19][2] = 8'h24;
frames[17][19][3] = 8'h48;
frames[17][19][4] = 8'h48;
frames[17][19][5] = 8'h48;
frames[17][19][6] = 8'h44;
frames[17][19][7] = 8'h24;
frames[17][19][8] = 8'h24;
frames[17][19][9] = 8'h24;
frames[17][19][10] = 8'h24;
frames[17][19][11] = 8'h24;
frames[17][19][12] = 8'h44;
frames[17][19][13] = 8'h44;
frames[17][19][14] = 8'h44;
frames[17][19][15] = 8'h44;
frames[17][19][16] = 8'h24;
frames[17][19][17] = 8'h24;
frames[17][19][18] = 8'h24;
frames[17][19][19] = 8'h24;
frames[17][19][20] = 8'h24;
frames[17][19][21] = 8'h24;
frames[17][19][22] = 8'h24;
frames[17][19][23] = 8'h24;
frames[17][19][24] = 8'h24;
frames[17][19][25] = 8'h24;
frames[17][19][26] = 8'h24;
frames[17][19][27] = 8'h00;
frames[17][19][28] = 8'h20;
frames[17][19][29] = 8'h24;
frames[17][19][30] = 8'h24;
frames[17][19][31] = 8'h24;
frames[17][19][32] = 8'h24;
frames[17][19][33] = 8'h24;
frames[17][19][34] = 8'h00;
frames[17][19][35] = 8'h00;
frames[17][19][36] = 8'h00;
frames[17][19][37] = 8'h00;
frames[17][19][38] = 8'h04;
frames[17][19][39] = 8'h04;
frames[17][20][0] = 8'h24;
frames[17][20][1] = 8'h24;
frames[17][20][2] = 8'h24;
frames[17][20][3] = 8'h24;
frames[17][20][4] = 8'h24;
frames[17][20][5] = 8'h44;
frames[17][20][6] = 8'h69;
frames[17][20][7] = 8'h48;
frames[17][20][8] = 8'h24;
frames[17][20][9] = 8'h24;
frames[17][20][10] = 8'h24;
frames[17][20][11] = 8'h24;
frames[17][20][12] = 8'h44;
frames[17][20][13] = 8'h44;
frames[17][20][14] = 8'h24;
frames[17][20][15] = 8'h24;
frames[17][20][16] = 8'h24;
frames[17][20][17] = 8'h24;
frames[17][20][18] = 8'h24;
frames[17][20][19] = 8'h24;
frames[17][20][20] = 8'h24;
frames[17][20][21] = 8'h24;
frames[17][20][22] = 8'h24;
frames[17][20][23] = 8'h24;
frames[17][20][24] = 8'h24;
frames[17][20][25] = 8'h24;
frames[17][20][26] = 8'h49;
frames[17][20][27] = 8'h4d;
frames[17][20][28] = 8'h49;
frames[17][20][29] = 8'h24;
frames[17][20][30] = 8'h04;
frames[17][20][31] = 8'h24;
frames[17][20][32] = 8'h24;
frames[17][20][33] = 8'h28;
frames[17][20][34] = 8'h24;
frames[17][20][35] = 8'h24;
frames[17][20][36] = 8'h28;
frames[17][20][37] = 8'h24;
frames[17][20][38] = 8'h00;
frames[17][20][39] = 8'h00;
frames[17][21][0] = 8'h24;
frames[17][21][1] = 8'h24;
frames[17][21][2] = 8'h04;
frames[17][21][3] = 8'h24;
frames[17][21][4] = 8'h24;
frames[17][21][5] = 8'h24;
frames[17][21][6] = 8'h24;
frames[17][21][7] = 8'h49;
frames[17][21][8] = 8'h49;
frames[17][21][9] = 8'h49;
frames[17][21][10] = 8'h44;
frames[17][21][11] = 8'h24;
frames[17][21][12] = 8'h24;
frames[17][21][13] = 8'h44;
frames[17][21][14] = 8'h24;
frames[17][21][15] = 8'h24;
frames[17][21][16] = 8'h24;
frames[17][21][17] = 8'h24;
frames[17][21][18] = 8'h24;
frames[17][21][19] = 8'h24;
frames[17][21][20] = 8'h24;
frames[17][21][21] = 8'h24;
frames[17][21][22] = 8'h24;
frames[17][21][23] = 8'h24;
frames[17][21][24] = 8'h24;
frames[17][21][25] = 8'h24;
frames[17][21][26] = 8'h6d;
frames[17][21][27] = 8'h71;
frames[17][21][28] = 8'h71;
frames[17][21][29] = 8'h6d;
frames[17][21][30] = 8'h24;
frames[17][21][31] = 8'h6d;
frames[17][21][32] = 8'h48;
frames[17][21][33] = 8'h4d;
frames[17][21][34] = 8'h24;
frames[17][21][35] = 8'h96;
frames[17][21][36] = 8'h92;
frames[17][21][37] = 8'h6d;
frames[17][21][38] = 8'h24;
frames[17][21][39] = 8'h00;
frames[17][22][0] = 8'h20;
frames[17][22][1] = 8'h24;
frames[17][22][2] = 8'h24;
frames[17][22][3] = 8'h24;
frames[17][22][4] = 8'h24;
frames[17][22][5] = 8'h24;
frames[17][22][6] = 8'h24;
frames[17][22][7] = 8'h24;
frames[17][22][8] = 8'h24;
frames[17][22][9] = 8'h49;
frames[17][22][10] = 8'h6d;
frames[17][22][11] = 8'h49;
frames[17][22][12] = 8'h44;
frames[17][22][13] = 8'h24;
frames[17][22][14] = 8'h44;
frames[17][22][15] = 8'h44;
frames[17][22][16] = 8'h44;
frames[17][22][17] = 8'h44;
frames[17][22][18] = 8'h44;
frames[17][22][19] = 8'h44;
frames[17][22][20] = 8'h44;
frames[17][22][21] = 8'h24;
frames[17][22][22] = 8'h24;
frames[17][22][23] = 8'h24;
frames[17][22][24] = 8'h24;
frames[17][22][25] = 8'h24;
frames[17][22][26] = 8'h4d;
frames[17][22][27] = 8'h71;
frames[17][22][28] = 8'h71;
frames[17][22][29] = 8'h4d;
frames[17][22][30] = 8'h24;
frames[17][22][31] = 8'h4d;
frames[17][22][32] = 8'h6d;
frames[17][22][33] = 8'h71;
frames[17][22][34] = 8'h49;
frames[17][22][35] = 8'h92;
frames[17][22][36] = 8'h92;
frames[17][22][37] = 8'h92;
frames[17][22][38] = 8'h24;
frames[17][22][39] = 8'h00;
frames[17][23][0] = 8'h20;
frames[17][23][1] = 8'h24;
frames[17][23][2] = 8'h24;
frames[17][23][3] = 8'h24;
frames[17][23][4] = 8'h24;
frames[17][23][5] = 8'h24;
frames[17][23][6] = 8'h24;
frames[17][23][7] = 8'h24;
frames[17][23][8] = 8'h24;
frames[17][23][9] = 8'h24;
frames[17][23][10] = 8'h44;
frames[17][23][11] = 8'h49;
frames[17][23][12] = 8'h6d;
frames[17][23][13] = 8'h49;
frames[17][23][14] = 8'h44;
frames[17][23][15] = 8'h44;
frames[17][23][16] = 8'h44;
frames[17][23][17] = 8'h44;
frames[17][23][18] = 8'h44;
frames[17][23][19] = 8'h44;
frames[17][23][20] = 8'h44;
frames[17][23][21] = 8'h24;
frames[17][23][22] = 8'h24;
frames[17][23][23] = 8'h44;
frames[17][23][24] = 8'h24;
frames[17][23][25] = 8'h24;
frames[17][23][26] = 8'h6d;
frames[17][23][27] = 8'h92;
frames[17][23][28] = 8'h71;
frames[17][23][29] = 8'h6d;
frames[17][23][30] = 8'h24;
frames[17][23][31] = 8'h24;
frames[17][23][32] = 8'h28;
frames[17][23][33] = 8'h6d;
frames[17][23][34] = 8'h49;
frames[17][23][35] = 8'h6d;
frames[17][23][36] = 8'h6e;
frames[17][23][37] = 8'h92;
frames[17][23][38] = 8'h24;
frames[17][23][39] = 8'h00;
frames[17][24][0] = 8'h00;
frames[17][24][1] = 8'h20;
frames[17][24][2] = 8'h24;
frames[17][24][3] = 8'h24;
frames[17][24][4] = 8'h24;
frames[17][24][5] = 8'h24;
frames[17][24][6] = 8'h24;
frames[17][24][7] = 8'h24;
frames[17][24][8] = 8'h24;
frames[17][24][9] = 8'h24;
frames[17][24][10] = 8'h24;
frames[17][24][11] = 8'h24;
frames[17][24][12] = 8'h48;
frames[17][24][13] = 8'h6d;
frames[17][24][14] = 8'h6d;
frames[17][24][15] = 8'h6d;
frames[17][24][16] = 8'h49;
frames[17][24][17] = 8'h48;
frames[17][24][18] = 8'h44;
frames[17][24][19] = 8'h44;
frames[17][24][20] = 8'h44;
frames[17][24][21] = 8'h24;
frames[17][24][22] = 8'h24;
frames[17][24][23] = 8'h48;
frames[17][24][24] = 8'h24;
frames[17][24][25] = 8'h24;
frames[17][24][26] = 8'h28;
frames[17][24][27] = 8'h24;
frames[17][24][28] = 8'h24;
frames[17][24][29] = 8'h48;
frames[17][24][30] = 8'h24;
frames[17][24][31] = 8'h24;
frames[17][24][32] = 8'h24;
frames[17][24][33] = 8'h24;
frames[17][24][34] = 8'h24;
frames[17][24][35] = 8'h24;
frames[17][24][36] = 8'h24;
frames[17][24][37] = 8'h25;
frames[17][24][38] = 8'h24;
frames[17][24][39] = 8'h24;
frames[17][25][0] = 8'h20;
frames[17][25][1] = 8'h20;
frames[17][25][2] = 8'h24;
frames[17][25][3] = 8'h24;
frames[17][25][4] = 8'h24;
frames[17][25][5] = 8'h24;
frames[17][25][6] = 8'h24;
frames[17][25][7] = 8'h24;
frames[17][25][8] = 8'h24;
frames[17][25][9] = 8'h24;
frames[17][25][10] = 8'h24;
frames[17][25][11] = 8'h24;
frames[17][25][12] = 8'h24;
frames[17][25][13] = 8'h24;
frames[17][25][14] = 8'h24;
frames[17][25][15] = 8'h6d;
frames[17][25][16] = 8'h6d;
frames[17][25][17] = 8'h49;
frames[17][25][18] = 8'h48;
frames[17][25][19] = 8'h44;
frames[17][25][20] = 8'h44;
frames[17][25][21] = 8'h24;
frames[17][25][22] = 8'h24;
frames[17][25][23] = 8'h24;
frames[17][25][24] = 8'h24;
frames[17][25][25] = 8'h24;
frames[17][25][26] = 8'h6d;
frames[17][25][27] = 8'h6d;
frames[17][25][28] = 8'h6d;
frames[17][25][29] = 8'h71;
frames[17][25][30] = 8'h6d;
frames[17][25][31] = 8'h6d;
frames[17][25][32] = 8'h6d;
frames[17][25][33] = 8'h49;
frames[17][25][34] = 8'h6d;
frames[17][25][35] = 8'h6d;
frames[17][25][36] = 8'h6d;
frames[17][25][37] = 8'h6d;
frames[17][25][38] = 8'h24;
frames[17][25][39] = 8'h24;
frames[17][26][0] = 8'h48;
frames[17][26][1] = 8'h00;
frames[17][26][2] = 8'h00;
frames[17][26][3] = 8'h24;
frames[17][26][4] = 8'h24;
frames[17][26][5] = 8'h24;
frames[17][26][6] = 8'h24;
frames[17][26][7] = 8'h24;
frames[17][26][8] = 8'h24;
frames[17][26][9] = 8'h24;
frames[17][26][10] = 8'h24;
frames[17][26][11] = 8'h24;
frames[17][26][12] = 8'h24;
frames[17][26][13] = 8'h24;
frames[17][26][14] = 8'h24;
frames[17][26][15] = 8'h24;
frames[17][26][16] = 8'h48;
frames[17][26][17] = 8'h6d;
frames[17][26][18] = 8'h6d;
frames[17][26][19] = 8'h49;
frames[17][26][20] = 8'h44;
frames[17][26][21] = 8'h24;
frames[17][26][22] = 8'h24;
frames[17][26][23] = 8'h24;
frames[17][26][24] = 8'h24;
frames[17][26][25] = 8'h24;
frames[17][26][26] = 8'h49;
frames[17][26][27] = 8'h6d;
frames[17][26][28] = 8'h91;
frames[17][26][29] = 8'h92;
frames[17][26][30] = 8'h92;
frames[17][26][31] = 8'h92;
frames[17][26][32] = 8'h6d;
frames[17][26][33] = 8'h24;
frames[17][26][34] = 8'h4d;
frames[17][26][35] = 8'h92;
frames[17][26][36] = 8'h6d;
frames[17][26][37] = 8'h49;
frames[17][26][38] = 8'h24;
frames[17][26][39] = 8'h04;
frames[17][27][0] = 8'h48;
frames[17][27][1] = 8'h00;
frames[17][27][2] = 8'h00;
frames[17][27][3] = 8'h04;
frames[17][27][4] = 8'h24;
frames[17][27][5] = 8'h24;
frames[17][27][6] = 8'h24;
frames[17][27][7] = 8'h24;
frames[17][27][8] = 8'h24;
frames[17][27][9] = 8'h24;
frames[17][27][10] = 8'h24;
frames[17][27][11] = 8'h24;
frames[17][27][12] = 8'h24;
frames[17][27][13] = 8'h24;
frames[17][27][14] = 8'h24;
frames[17][27][15] = 8'h24;
frames[17][27][16] = 8'h24;
frames[17][27][17] = 8'h24;
frames[17][27][18] = 8'h48;
frames[17][27][19] = 8'h6d;
frames[17][27][20] = 8'h6d;
frames[17][27][21] = 8'h48;
frames[17][27][22] = 8'h24;
frames[17][27][23] = 8'h24;
frames[17][27][24] = 8'h24;
frames[17][27][25] = 8'h24;
frames[17][27][26] = 8'h49;
frames[17][27][27] = 8'h6d;
frames[17][27][28] = 8'h92;
frames[17][27][29] = 8'h91;
frames[17][27][30] = 8'h92;
frames[17][27][31] = 8'h92;
frames[17][27][32] = 8'h92;
frames[17][27][33] = 8'h49;
frames[17][27][34] = 8'h6d;
frames[17][27][35] = 8'h92;
frames[17][27][36] = 8'h91;
frames[17][27][37] = 8'h6d;
frames[17][27][38] = 8'h24;
frames[17][27][39] = 8'h04;
frames[17][28][0] = 8'h6d;
frames[17][28][1] = 8'h20;
frames[17][28][2] = 8'h00;
frames[17][28][3] = 8'h00;
frames[17][28][4] = 8'h24;
frames[17][28][5] = 8'h24;
frames[17][28][6] = 8'h24;
frames[17][28][7] = 8'h24;
frames[17][28][8] = 8'h24;
frames[17][28][9] = 8'h24;
frames[17][28][10] = 8'h24;
frames[17][28][11] = 8'h24;
frames[17][28][12] = 8'h24;
frames[17][28][13] = 8'h24;
frames[17][28][14] = 8'h24;
frames[17][28][15] = 8'h24;
frames[17][28][16] = 8'h24;
frames[17][28][17] = 8'h24;
frames[17][28][18] = 8'h24;
frames[17][28][19] = 8'h24;
frames[17][28][20] = 8'h48;
frames[17][28][21] = 8'h49;
frames[17][28][22] = 8'h6d;
frames[17][28][23] = 8'h49;
frames[17][28][24] = 8'h24;
frames[17][28][25] = 8'h24;
frames[17][28][26] = 8'h24;
frames[17][28][27] = 8'h49;
frames[17][28][28] = 8'h49;
frames[17][28][29] = 8'h49;
frames[17][28][30] = 8'h49;
frames[17][28][31] = 8'h49;
frames[17][28][32] = 8'h49;
frames[17][28][33] = 8'h24;
frames[17][28][34] = 8'h49;
frames[17][28][35] = 8'h49;
frames[17][28][36] = 8'h49;
frames[17][28][37] = 8'h4d;
frames[17][28][38] = 8'h24;
frames[17][28][39] = 8'h00;
frames[17][29][0] = 8'h92;
frames[17][29][1] = 8'h92;
frames[17][29][2] = 8'h24;
frames[17][29][3] = 8'h24;
frames[17][29][4] = 8'h24;
frames[17][29][5] = 8'h24;
frames[17][29][6] = 8'h24;
frames[17][29][7] = 8'h24;
frames[17][29][8] = 8'h24;
frames[17][29][9] = 8'h24;
frames[17][29][10] = 8'h24;
frames[17][29][11] = 8'h24;
frames[17][29][12] = 8'h24;
frames[17][29][13] = 8'h24;
frames[17][29][14] = 8'h24;
frames[17][29][15] = 8'h24;
frames[17][29][16] = 8'h24;
frames[17][29][17] = 8'h24;
frames[17][29][18] = 8'h24;
frames[17][29][19] = 8'h24;
frames[17][29][20] = 8'h24;
frames[17][29][21] = 8'h24;
frames[17][29][22] = 8'h44;
frames[17][29][23] = 8'h69;
frames[17][29][24] = 8'h49;
frames[17][29][25] = 8'h44;
frames[17][29][26] = 8'h24;
frames[17][29][27] = 8'h00;
frames[17][29][28] = 8'h00;
frames[17][29][29] = 8'h04;
frames[17][29][30] = 8'h04;
frames[17][29][31] = 8'h04;
frames[17][29][32] = 8'h00;
frames[17][29][33] = 8'h24;
frames[17][29][34] = 8'h00;
frames[17][29][35] = 8'h00;
frames[17][29][36] = 8'h00;
frames[17][29][37] = 8'h00;
frames[17][29][38] = 8'h00;
frames[17][29][39] = 8'h04;
frames[18][0][0] = 8'hf6;
frames[18][0][1] = 8'hfa;
frames[18][0][2] = 8'hd6;
frames[18][0][3] = 8'hd6;
frames[18][0][4] = 8'hd6;
frames[18][0][5] = 8'hfa;
frames[18][0][6] = 8'h6d;
frames[18][0][7] = 8'h44;
frames[18][0][8] = 8'h48;
frames[18][0][9] = 8'h48;
frames[18][0][10] = 8'h48;
frames[18][0][11] = 8'h44;
frames[18][0][12] = 8'h44;
frames[18][0][13] = 8'h48;
frames[18][0][14] = 8'h44;
frames[18][0][15] = 8'h44;
frames[18][0][16] = 8'h48;
frames[18][0][17] = 8'h44;
frames[18][0][18] = 8'h24;
frames[18][0][19] = 8'h48;
frames[18][0][20] = 8'h48;
frames[18][0][21] = 8'h44;
frames[18][0][22] = 8'h44;
frames[18][0][23] = 8'h48;
frames[18][0][24] = 8'h49;
frames[18][0][25] = 8'h44;
frames[18][0][26] = 8'h44;
frames[18][0][27] = 8'h49;
frames[18][0][28] = 8'h49;
frames[18][0][29] = 8'h48;
frames[18][0][30] = 8'h24;
frames[18][0][31] = 8'h44;
frames[18][0][32] = 8'h44;
frames[18][0][33] = 8'h24;
frames[18][0][34] = 8'h44;
frames[18][0][35] = 8'h24;
frames[18][0][36] = 8'h00;
frames[18][0][37] = 8'h48;
frames[18][0][38] = 8'h24;
frames[18][0][39] = 8'h00;
frames[18][1][0] = 8'hd6;
frames[18][1][1] = 8'hf6;
frames[18][1][2] = 8'hfa;
frames[18][1][3] = 8'hfa;
frames[18][1][4] = 8'hf6;
frames[18][1][5] = 8'hfa;
frames[18][1][6] = 8'hfa;
frames[18][1][7] = 8'h69;
frames[18][1][8] = 8'h44;
frames[18][1][9] = 8'h48;
frames[18][1][10] = 8'h44;
frames[18][1][11] = 8'h44;
frames[18][1][12] = 8'h44;
frames[18][1][13] = 8'h48;
frames[18][1][14] = 8'h44;
frames[18][1][15] = 8'h44;
frames[18][1][16] = 8'h48;
frames[18][1][17] = 8'h44;
frames[18][1][18] = 8'h44;
frames[18][1][19] = 8'h48;
frames[18][1][20] = 8'h48;
frames[18][1][21] = 8'h44;
frames[18][1][22] = 8'h44;
frames[18][1][23] = 8'h69;
frames[18][1][24] = 8'h48;
frames[18][1][25] = 8'h44;
frames[18][1][26] = 8'h44;
frames[18][1][27] = 8'h49;
frames[18][1][28] = 8'h69;
frames[18][1][29] = 8'h48;
frames[18][1][30] = 8'h44;
frames[18][1][31] = 8'h48;
frames[18][1][32] = 8'h44;
frames[18][1][33] = 8'h44;
frames[18][1][34] = 8'h44;
frames[18][1][35] = 8'h24;
frames[18][1][36] = 8'h49;
frames[18][1][37] = 8'hb6;
frames[18][1][38] = 8'hb6;
frames[18][1][39] = 8'h24;
frames[18][2][0] = 8'hd6;
frames[18][2][1] = 8'hd6;
frames[18][2][2] = 8'hf6;
frames[18][2][3] = 8'hfa;
frames[18][2][4] = 8'hfa;
frames[18][2][5] = 8'hfa;
frames[18][2][6] = 8'hfa;
frames[18][2][7] = 8'hf6;
frames[18][2][8] = 8'h8d;
frames[18][2][9] = 8'h68;
frames[18][2][10] = 8'h44;
frames[18][2][11] = 8'h44;
frames[18][2][12] = 8'h44;
frames[18][2][13] = 8'h48;
frames[18][2][14] = 8'h44;
frames[18][2][15] = 8'h44;
frames[18][2][16] = 8'h48;
frames[18][2][17] = 8'h48;
frames[18][2][18] = 8'h44;
frames[18][2][19] = 8'h44;
frames[18][2][20] = 8'h48;
frames[18][2][21] = 8'h44;
frames[18][2][22] = 8'h44;
frames[18][2][23] = 8'h69;
frames[18][2][24] = 8'h49;
frames[18][2][25] = 8'h48;
frames[18][2][26] = 8'h48;
frames[18][2][27] = 8'h69;
frames[18][2][28] = 8'h69;
frames[18][2][29] = 8'h48;
frames[18][2][30] = 8'h48;
frames[18][2][31] = 8'h48;
frames[18][2][32] = 8'h44;
frames[18][2][33] = 8'h48;
frames[18][2][34] = 8'h44;
frames[18][2][35] = 8'h24;
frames[18][2][36] = 8'h92;
frames[18][2][37] = 8'h6d;
frames[18][2][38] = 8'h4d;
frames[18][2][39] = 8'h4e;
frames[18][3][0] = 8'hd6;
frames[18][3][1] = 8'hd6;
frames[18][3][2] = 8'hd6;
frames[18][3][3] = 8'hd6;
frames[18][3][4] = 8'hf6;
frames[18][3][5] = 8'hf6;
frames[18][3][6] = 8'hf6;
frames[18][3][7] = 8'hf6;
frames[18][3][8] = 8'hfa;
frames[18][3][9] = 8'hd6;
frames[18][3][10] = 8'h6d;
frames[18][3][11] = 8'h44;
frames[18][3][12] = 8'h44;
frames[18][3][13] = 8'h48;
frames[18][3][14] = 8'h44;
frames[18][3][15] = 8'h44;
frames[18][3][16] = 8'h48;
frames[18][3][17] = 8'h48;
frames[18][3][18] = 8'h44;
frames[18][3][19] = 8'h48;
frames[18][3][20] = 8'h48;
frames[18][3][21] = 8'h48;
frames[18][3][22] = 8'h48;
frames[18][3][23] = 8'h69;
frames[18][3][24] = 8'h69;
frames[18][3][25] = 8'h49;
frames[18][3][26] = 8'h48;
frames[18][3][27] = 8'h44;
frames[18][3][28] = 8'h24;
frames[18][3][29] = 8'h44;
frames[18][3][30] = 8'h24;
frames[18][3][31] = 8'h24;
frames[18][3][32] = 8'h24;
frames[18][3][33] = 8'h24;
frames[18][3][34] = 8'h24;
frames[18][3][35] = 8'h48;
frames[18][3][36] = 8'h92;
frames[18][3][37] = 8'h92;
frames[18][3][38] = 8'h49;
frames[18][3][39] = 8'h72;
frames[18][4][0] = 8'hb1;
frames[18][4][1] = 8'hd2;
frames[18][4][2] = 8'hd2;
frames[18][4][3] = 8'hd6;
frames[18][4][4] = 8'hd6;
frames[18][4][5] = 8'hd6;
frames[18][4][6] = 8'hd6;
frames[18][4][7] = 8'hf6;
frames[18][4][8] = 8'hf6;
frames[18][4][9] = 8'hfa;
frames[18][4][10] = 8'hfa;
frames[18][4][11] = 8'hb1;
frames[18][4][12] = 8'h68;
frames[18][4][13] = 8'h48;
frames[18][4][14] = 8'h44;
frames[18][4][15] = 8'h69;
frames[18][4][16] = 8'h68;
frames[18][4][17] = 8'h48;
frames[18][4][18] = 8'h49;
frames[18][4][19] = 8'h48;
frames[18][4][20] = 8'h48;
frames[18][4][21] = 8'h48;
frames[18][4][22] = 8'h48;
frames[18][4][23] = 8'h44;
frames[18][4][24] = 8'h44;
frames[18][4][25] = 8'h44;
frames[18][4][26] = 8'h24;
frames[18][4][27] = 8'h24;
frames[18][4][28] = 8'h24;
frames[18][4][29] = 8'h24;
frames[18][4][30] = 8'h24;
frames[18][4][31] = 8'h24;
frames[18][4][32] = 8'h24;
frames[18][4][33] = 8'h24;
frames[18][4][34] = 8'h24;
frames[18][4][35] = 8'h24;
frames[18][4][36] = 8'h92;
frames[18][4][37] = 8'h6d;
frames[18][4][38] = 8'h6e;
frames[18][4][39] = 8'h6e;
frames[18][5][0] = 8'had;
frames[18][5][1] = 8'hb1;
frames[18][5][2] = 8'hd1;
frames[18][5][3] = 8'hd2;
frames[18][5][4] = 8'hd2;
frames[18][5][5] = 8'hd2;
frames[18][5][6] = 8'hd2;
frames[18][5][7] = 8'hd6;
frames[18][5][8] = 8'hd6;
frames[18][5][9] = 8'hf6;
frames[18][5][10] = 8'hf6;
frames[18][5][11] = 8'hfa;
frames[18][5][12] = 8'hf6;
frames[18][5][13] = 8'hb2;
frames[18][5][14] = 8'h69;
frames[18][5][15] = 8'h44;
frames[18][5][16] = 8'h44;
frames[18][5][17] = 8'h48;
frames[18][5][18] = 8'h48;
frames[18][5][19] = 8'h44;
frames[18][5][20] = 8'h44;
frames[18][5][21] = 8'h48;
frames[18][5][22] = 8'h44;
frames[18][5][23] = 8'h44;
frames[18][5][24] = 8'h24;
frames[18][5][25] = 8'h24;
frames[18][5][26] = 8'h24;
frames[18][5][27] = 8'h24;
frames[18][5][28] = 8'h24;
frames[18][5][29] = 8'h24;
frames[18][5][30] = 8'h24;
frames[18][5][31] = 8'h24;
frames[18][5][32] = 8'h24;
frames[18][5][33] = 8'h24;
frames[18][5][34] = 8'h24;
frames[18][5][35] = 8'h24;
frames[18][5][36] = 8'h49;
frames[18][5][37] = 8'h92;
frames[18][5][38] = 8'h92;
frames[18][5][39] = 8'h24;
frames[18][6][0] = 8'h8d;
frames[18][6][1] = 8'h8d;
frames[18][6][2] = 8'had;
frames[18][6][3] = 8'hb1;
frames[18][6][4] = 8'hb1;
frames[18][6][5] = 8'hb1;
frames[18][6][6] = 8'hd2;
frames[18][6][7] = 8'hd2;
frames[18][6][8] = 8'hd2;
frames[18][6][9] = 8'hd6;
frames[18][6][10] = 8'hf6;
frames[18][6][11] = 8'hf6;
frames[18][6][12] = 8'hf6;
frames[18][6][13] = 8'hfa;
frames[18][6][14] = 8'hfa;
frames[18][6][15] = 8'h8d;
frames[18][6][16] = 8'h44;
frames[18][6][17] = 8'h48;
frames[18][6][18] = 8'h48;
frames[18][6][19] = 8'h44;
frames[18][6][20] = 8'h44;
frames[18][6][21] = 8'h44;
frames[18][6][22] = 8'h44;
frames[18][6][23] = 8'h44;
frames[18][6][24] = 8'h24;
frames[18][6][25] = 8'h24;
frames[18][6][26] = 8'h24;
frames[18][6][27] = 8'h24;
frames[18][6][28] = 8'h24;
frames[18][6][29] = 8'h24;
frames[18][6][30] = 8'h24;
frames[18][6][31] = 8'h24;
frames[18][6][32] = 8'h24;
frames[18][6][33] = 8'h24;
frames[18][6][34] = 8'h24;
frames[18][6][35] = 8'h24;
frames[18][6][36] = 8'h24;
frames[18][6][37] = 8'h24;
frames[18][6][38] = 8'h24;
frames[18][6][39] = 8'h24;
frames[18][7][0] = 8'h69;
frames[18][7][1] = 8'h89;
frames[18][7][2] = 8'h8d;
frames[18][7][3] = 8'had;
frames[18][7][4] = 8'hb1;
frames[18][7][5] = 8'hb1;
frames[18][7][6] = 8'hd2;
frames[18][7][7] = 8'hd2;
frames[18][7][8] = 8'hd2;
frames[18][7][9] = 8'hd2;
frames[18][7][10] = 8'hd6;
frames[18][7][11] = 8'hf6;
frames[18][7][12] = 8'hf6;
frames[18][7][13] = 8'hfa;
frames[18][7][14] = 8'hfa;
frames[18][7][15] = 8'hf6;
frames[18][7][16] = 8'h6d;
frames[18][7][17] = 8'h44;
frames[18][7][18] = 8'h48;
frames[18][7][19] = 8'h48;
frames[18][7][20] = 8'h44;
frames[18][7][21] = 8'h44;
frames[18][7][22] = 8'h44;
frames[18][7][23] = 8'h44;
frames[18][7][24] = 8'h24;
frames[18][7][25] = 8'h24;
frames[18][7][26] = 8'h24;
frames[18][7][27] = 8'h24;
frames[18][7][28] = 8'h24;
frames[18][7][29] = 8'h24;
frames[18][7][30] = 8'h24;
frames[18][7][31] = 8'h24;
frames[18][7][32] = 8'h24;
frames[18][7][33] = 8'h24;
frames[18][7][34] = 8'h24;
frames[18][7][35] = 8'h24;
frames[18][7][36] = 8'h24;
frames[18][7][37] = 8'h24;
frames[18][7][38] = 8'h24;
frames[18][7][39] = 8'h24;
frames[18][8][0] = 8'h68;
frames[18][8][1] = 8'h68;
frames[18][8][2] = 8'h68;
frames[18][8][3] = 8'h8d;
frames[18][8][4] = 8'h8d;
frames[18][8][5] = 8'had;
frames[18][8][6] = 8'hb1;
frames[18][8][7] = 8'hb1;
frames[18][8][8] = 8'hd1;
frames[18][8][9] = 8'hd1;
frames[18][8][10] = 8'hd2;
frames[18][8][11] = 8'hd6;
frames[18][8][12] = 8'hf6;
frames[18][8][13] = 8'hfa;
frames[18][8][14] = 8'hfa;
frames[18][8][15] = 8'hfa;
frames[18][8][16] = 8'hfa;
frames[18][8][17] = 8'h8d;
frames[18][8][18] = 8'h48;
frames[18][8][19] = 8'h44;
frames[18][8][20] = 8'h44;
frames[18][8][21] = 8'h44;
frames[18][8][22] = 8'h24;
frames[18][8][23] = 8'h24;
frames[18][8][24] = 8'h24;
frames[18][8][25] = 8'h24;
frames[18][8][26] = 8'h24;
frames[18][8][27] = 8'h24;
frames[18][8][28] = 8'h24;
frames[18][8][29] = 8'h24;
frames[18][8][30] = 8'h24;
frames[18][8][31] = 8'h24;
frames[18][8][32] = 8'h24;
frames[18][8][33] = 8'h24;
frames[18][8][34] = 8'h24;
frames[18][8][35] = 8'h24;
frames[18][8][36] = 8'h24;
frames[18][8][37] = 8'h24;
frames[18][8][38] = 8'h24;
frames[18][8][39] = 8'h24;
frames[18][9][0] = 8'h48;
frames[18][9][1] = 8'h48;
frames[18][9][2] = 8'h68;
frames[18][9][3] = 8'h68;
frames[18][9][4] = 8'h69;
frames[18][9][5] = 8'h8d;
frames[18][9][6] = 8'had;
frames[18][9][7] = 8'hb1;
frames[18][9][8] = 8'hb1;
frames[18][9][9] = 8'hb1;
frames[18][9][10] = 8'hd1;
frames[18][9][11] = 8'hd2;
frames[18][9][12] = 8'hd6;
frames[18][9][13] = 8'hf6;
frames[18][9][14] = 8'hf6;
frames[18][9][15] = 8'hfa;
frames[18][9][16] = 8'hfa;
frames[18][9][17] = 8'hfa;
frames[18][9][18] = 8'hd6;
frames[18][9][19] = 8'h69;
frames[18][9][20] = 8'h24;
frames[18][9][21] = 8'h24;
frames[18][9][22] = 8'h24;
frames[18][9][23] = 8'h24;
frames[18][9][24] = 8'h24;
frames[18][9][25] = 8'h24;
frames[18][9][26] = 8'h24;
frames[18][9][27] = 8'h24;
frames[18][9][28] = 8'h24;
frames[18][9][29] = 8'h24;
frames[18][9][30] = 8'h24;
frames[18][9][31] = 8'h24;
frames[18][9][32] = 8'h24;
frames[18][9][33] = 8'h24;
frames[18][9][34] = 8'h24;
frames[18][9][35] = 8'h24;
frames[18][9][36] = 8'h24;
frames[18][9][37] = 8'h24;
frames[18][9][38] = 8'h24;
frames[18][9][39] = 8'h24;
frames[18][10][0] = 8'h6d;
frames[18][10][1] = 8'h91;
frames[18][10][2] = 8'h8d;
frames[18][10][3] = 8'h69;
frames[18][10][4] = 8'h69;
frames[18][10][5] = 8'h69;
frames[18][10][6] = 8'h69;
frames[18][10][7] = 8'h89;
frames[18][10][8] = 8'h8d;
frames[18][10][9] = 8'had;
frames[18][10][10] = 8'hb1;
frames[18][10][11] = 8'hb1;
frames[18][10][12] = 8'hd2;
frames[18][10][13] = 8'hd6;
frames[18][10][14] = 8'hd6;
frames[18][10][15] = 8'hf6;
frames[18][10][16] = 8'hf6;
frames[18][10][17] = 8'hfa;
frames[18][10][18] = 8'hfa;
frames[18][10][19] = 8'hfa;
frames[18][10][20] = 8'hb2;
frames[18][10][21] = 8'h68;
frames[18][10][22] = 8'h24;
frames[18][10][23] = 8'h24;
frames[18][10][24] = 8'h24;
frames[18][10][25] = 8'h24;
frames[18][10][26] = 8'h24;
frames[18][10][27] = 8'h44;
frames[18][10][28] = 8'h6d;
frames[18][10][29] = 8'hb6;
frames[18][10][30] = 8'hda;
frames[18][10][31] = 8'hda;
frames[18][10][32] = 8'hda;
frames[18][10][33] = 8'h92;
frames[18][10][34] = 8'h49;
frames[18][10][35] = 8'h24;
frames[18][10][36] = 8'h24;
frames[18][10][37] = 8'h24;
frames[18][10][38] = 8'h24;
frames[18][10][39] = 8'h24;
frames[18][11][0] = 8'hda;
frames[18][11][1] = 8'hda;
frames[18][11][2] = 8'hb6;
frames[18][11][3] = 8'hb6;
frames[18][11][4] = 8'h92;
frames[18][11][5] = 8'h92;
frames[18][11][6] = 8'h91;
frames[18][11][7] = 8'h8d;
frames[18][11][8] = 8'h69;
frames[18][11][9] = 8'h69;
frames[18][11][10] = 8'h8d;
frames[18][11][11] = 8'hb1;
frames[18][11][12] = 8'hd1;
frames[18][11][13] = 8'hd2;
frames[18][11][14] = 8'hd6;
frames[18][11][15] = 8'hf6;
frames[18][11][16] = 8'hf6;
frames[18][11][17] = 8'hf6;
frames[18][11][18] = 8'hf6;
frames[18][11][19] = 8'hf6;
frames[18][11][20] = 8'hfa;
frames[18][11][21] = 8'hd6;
frames[18][11][22] = 8'h48;
frames[18][11][23] = 8'h24;
frames[18][11][24] = 8'h48;
frames[18][11][25] = 8'h6d;
frames[18][11][26] = 8'hb2;
frames[18][11][27] = 8'hdb;
frames[18][11][28] = 8'hff;
frames[18][11][29] = 8'hff;
frames[18][11][30] = 8'hff;
frames[18][11][31] = 8'hff;
frames[18][11][32] = 8'hff;
frames[18][11][33] = 8'hff;
frames[18][11][34] = 8'hff;
frames[18][11][35] = 8'hb6;
frames[18][11][36] = 8'h49;
frames[18][11][37] = 8'h24;
frames[18][11][38] = 8'h24;
frames[18][11][39] = 8'h24;
frames[18][12][0] = 8'hb6;
frames[18][12][1] = 8'hb6;
frames[18][12][2] = 8'hba;
frames[18][12][3] = 8'hdb;
frames[18][12][4] = 8'hdb;
frames[18][12][5] = 8'hdf;
frames[18][12][6] = 8'hff;
frames[18][12][7] = 8'hff;
frames[18][12][8] = 8'hda;
frames[18][12][9] = 8'h44;
frames[18][12][10] = 8'h68;
frames[18][12][11] = 8'h8d;
frames[18][12][12] = 8'hb1;
frames[18][12][13] = 8'hd2;
frames[18][12][14] = 8'hd6;
frames[18][12][15] = 8'hf6;
frames[18][12][16] = 8'hf6;
frames[18][12][17] = 8'hf6;
frames[18][12][18] = 8'hf6;
frames[18][12][19] = 8'hf6;
frames[18][12][20] = 8'hf6;
frames[18][12][21] = 8'hd6;
frames[18][12][22] = 8'h91;
frames[18][12][23] = 8'hb6;
frames[18][12][24] = 8'hff;
frames[18][12][25] = 8'hff;
frames[18][12][26] = 8'hff;
frames[18][12][27] = 8'hff;
frames[18][12][28] = 8'hff;
frames[18][12][29] = 8'hff;
frames[18][12][30] = 8'hff;
frames[18][12][31] = 8'hff;
frames[18][12][32] = 8'hff;
frames[18][12][33] = 8'hff;
frames[18][12][34] = 8'hff;
frames[18][12][35] = 8'hff;
frames[18][12][36] = 8'hff;
frames[18][12][37] = 8'h91;
frames[18][12][38] = 8'h20;
frames[18][12][39] = 8'h24;
frames[18][13][0] = 8'hdb;
frames[18][13][1] = 8'hdf;
frames[18][13][2] = 8'hdf;
frames[18][13][3] = 8'hdf;
frames[18][13][4] = 8'hff;
frames[18][13][5] = 8'hff;
frames[18][13][6] = 8'hff;
frames[18][13][7] = 8'hff;
frames[18][13][8] = 8'h92;
frames[18][13][9] = 8'h00;
frames[18][13][10] = 8'h68;
frames[18][13][11] = 8'h8d;
frames[18][13][12] = 8'had;
frames[18][13][13] = 8'hb1;
frames[18][13][14] = 8'hd2;
frames[18][13][15] = 8'hd6;
frames[18][13][16] = 8'hd6;
frames[18][13][17] = 8'hf6;
frames[18][13][18] = 8'hd6;
frames[18][13][19] = 8'hf6;
frames[18][13][20] = 8'hf6;
frames[18][13][21] = 8'had;
frames[18][13][22] = 8'hb2;
frames[18][13][23] = 8'hff;
frames[18][13][24] = 8'hff;
frames[18][13][25] = 8'hff;
frames[18][13][26] = 8'hff;
frames[18][13][27] = 8'hff;
frames[18][13][28] = 8'hff;
frames[18][13][29] = 8'hff;
frames[18][13][30] = 8'hff;
frames[18][13][31] = 8'hff;
frames[18][13][32] = 8'hff;
frames[18][13][33] = 8'hff;
frames[18][13][34] = 8'hff;
frames[18][13][35] = 8'hff;
frames[18][13][36] = 8'hff;
frames[18][13][37] = 8'hff;
frames[18][13][38] = 8'h6d;
frames[18][13][39] = 8'h00;
frames[18][14][0] = 8'hdb;
frames[18][14][1] = 8'hdb;
frames[18][14][2] = 8'hdf;
frames[18][14][3] = 8'hdf;
frames[18][14][4] = 8'hff;
frames[18][14][5] = 8'hff;
frames[18][14][6] = 8'hff;
frames[18][14][7] = 8'hdb;
frames[18][14][8] = 8'h6d;
frames[18][14][9] = 8'h91;
frames[18][14][10] = 8'hfb;
frames[18][14][11] = 8'hda;
frames[18][14][12] = 8'h8d;
frames[18][14][13] = 8'had;
frames[18][14][14] = 8'hb1;
frames[18][14][15] = 8'hd2;
frames[18][14][16] = 8'hd2;
frames[18][14][17] = 8'hd6;
frames[18][14][18] = 8'hf6;
frames[18][14][19] = 8'hb2;
frames[18][14][20] = 8'hb1;
frames[18][14][21] = 8'h89;
frames[18][14][22] = 8'h8d;
frames[18][14][23] = 8'hff;
frames[18][14][24] = 8'hff;
frames[18][14][25] = 8'hff;
frames[18][14][26] = 8'hff;
frames[18][14][27] = 8'hff;
frames[18][14][28] = 8'hff;
frames[18][14][29] = 8'hff;
frames[18][14][30] = 8'hff;
frames[18][14][31] = 8'hff;
frames[18][14][32] = 8'hff;
frames[18][14][33] = 8'hff;
frames[18][14][34] = 8'hff;
frames[18][14][35] = 8'hff;
frames[18][14][36] = 8'hff;
frames[18][14][37] = 8'hff;
frames[18][14][38] = 8'hdb;
frames[18][14][39] = 8'h24;
frames[18][15][0] = 8'hdb;
frames[18][15][1] = 8'hdb;
frames[18][15][2] = 8'hba;
frames[18][15][3] = 8'h96;
frames[18][15][4] = 8'h71;
frames[18][15][5] = 8'h6d;
frames[18][15][6] = 8'h49;
frames[18][15][7] = 8'h6d;
frames[18][15][8] = 8'hfb;
frames[18][15][9] = 8'hff;
frames[18][15][10] = 8'hff;
frames[18][15][11] = 8'hff;
frames[18][15][12] = 8'hd6;
frames[18][15][13] = 8'h8d;
frames[18][15][14] = 8'had;
frames[18][15][15] = 8'hb1;
frames[18][15][16] = 8'hd1;
frames[18][15][17] = 8'hd2;
frames[18][15][18] = 8'hd6;
frames[18][15][19] = 8'h8d;
frames[18][15][20] = 8'h64;
frames[18][15][21] = 8'h69;
frames[18][15][22] = 8'h68;
frames[18][15][23] = 8'hd6;
frames[18][15][24] = 8'hfa;
frames[18][15][25] = 8'hff;
frames[18][15][26] = 8'hff;
frames[18][15][27] = 8'hff;
frames[18][15][28] = 8'hff;
frames[18][15][29] = 8'hff;
frames[18][15][30] = 8'hff;
frames[18][15][31] = 8'hff;
frames[18][15][32] = 8'hff;
frames[18][15][33] = 8'hff;
frames[18][15][34] = 8'hff;
frames[18][15][35] = 8'hff;
frames[18][15][36] = 8'hff;
frames[18][15][37] = 8'hff;
frames[18][15][38] = 8'hb6;
frames[18][15][39] = 8'h24;
frames[18][16][0] = 8'h69;
frames[18][16][1] = 8'h44;
frames[18][16][2] = 8'h24;
frames[18][16][3] = 8'h24;
frames[18][16][4] = 8'h24;
frames[18][16][5] = 8'h04;
frames[18][16][6] = 8'h20;
frames[18][16][7] = 8'hd6;
frames[18][16][8] = 8'hff;
frames[18][16][9] = 8'hff;
frames[18][16][10] = 8'hff;
frames[18][16][11] = 8'hff;
frames[18][16][12] = 8'hff;
frames[18][16][13] = 8'hb6;
frames[18][16][14] = 8'h89;
frames[18][16][15] = 8'had;
frames[18][16][16] = 8'hd1;
frames[18][16][17] = 8'hb1;
frames[18][16][18] = 8'h8d;
frames[18][16][19] = 8'h68;
frames[18][16][20] = 8'h44;
frames[18][16][21] = 8'h69;
frames[18][16][22] = 8'h68;
frames[18][16][23] = 8'h8d;
frames[18][16][24] = 8'hd6;
frames[18][16][25] = 8'hff;
frames[18][16][26] = 8'hff;
frames[18][16][27] = 8'hff;
frames[18][16][28] = 8'hff;
frames[18][16][29] = 8'hff;
frames[18][16][30] = 8'hff;
frames[18][16][31] = 8'hff;
frames[18][16][32] = 8'hff;
frames[18][16][33] = 8'hff;
frames[18][16][34] = 8'hff;
frames[18][16][35] = 8'hff;
frames[18][16][36] = 8'hda;
frames[18][16][37] = 8'hd6;
frames[18][16][38] = 8'h49;
frames[18][16][39] = 8'h00;
frames[18][17][0] = 8'h44;
frames[18][17][1] = 8'h24;
frames[18][17][2] = 8'h24;
frames[18][17][3] = 8'h24;
frames[18][17][4] = 8'h24;
frames[18][17][5] = 8'h00;
frames[18][17][6] = 8'h24;
frames[18][17][7] = 8'hfb;
frames[18][17][8] = 8'hff;
frames[18][17][9] = 8'hff;
frames[18][17][10] = 8'hff;
frames[18][17][11] = 8'hff;
frames[18][17][12] = 8'hff;
frames[18][17][13] = 8'hff;
frames[18][17][14] = 8'hd6;
frames[18][17][15] = 8'h8d;
frames[18][17][16] = 8'had;
frames[18][17][17] = 8'h8d;
frames[18][17][18] = 8'h64;
frames[18][17][19] = 8'h68;
frames[18][17][20] = 8'h44;
frames[18][17][21] = 8'h68;
frames[18][17][22] = 8'h68;
frames[18][17][23] = 8'h69;
frames[18][17][24] = 8'hd6;
frames[18][17][25] = 8'hff;
frames[18][17][26] = 8'hff;
frames[18][17][27] = 8'hff;
frames[18][17][28] = 8'hff;
frames[18][17][29] = 8'hfb;
frames[18][17][30] = 8'hfa;
frames[18][17][31] = 8'hda;
frames[18][17][32] = 8'hd6;
frames[18][17][33] = 8'hb6;
frames[18][17][34] = 8'hb1;
frames[18][17][35] = 8'h8d;
frames[18][17][36] = 8'h64;
frames[18][17][37] = 8'h68;
frames[18][17][38] = 8'h24;
frames[18][17][39] = 8'h00;
frames[18][18][0] = 8'h24;
frames[18][18][1] = 8'h49;
frames[18][18][2] = 8'h49;
frames[18][18][3] = 8'h24;
frames[18][18][4] = 8'h24;
frames[18][18][5] = 8'h24;
frames[18][18][6] = 8'h24;
frames[18][18][7] = 8'hfb;
frames[18][18][8] = 8'hff;
frames[18][18][9] = 8'hff;
frames[18][18][10] = 8'hff;
frames[18][18][11] = 8'hff;
frames[18][18][12] = 8'hff;
frames[18][18][13] = 8'hff;
frames[18][18][14] = 8'hff;
frames[18][18][15] = 8'hb1;
frames[18][18][16] = 8'h44;
frames[18][18][17] = 8'h44;
frames[18][18][18] = 8'h44;
frames[18][18][19] = 8'h68;
frames[18][18][20] = 8'h68;
frames[18][18][21] = 8'h44;
frames[18][18][22] = 8'h48;
frames[18][18][23] = 8'h44;
frames[18][18][24] = 8'h48;
frames[18][18][25] = 8'h6d;
frames[18][18][26] = 8'h8d;
frames[18][18][27] = 8'h8d;
frames[18][18][28] = 8'hb1;
frames[18][18][29] = 8'had;
frames[18][18][30] = 8'h8d;
frames[18][18][31] = 8'h8d;
frames[18][18][32] = 8'hb1;
frames[18][18][33] = 8'hb1;
frames[18][18][34] = 8'hb1;
frames[18][18][35] = 8'h8d;
frames[18][18][36] = 8'h44;
frames[18][18][37] = 8'h24;
frames[18][18][38] = 8'h00;
frames[18][18][39] = 8'h20;
frames[18][19][0] = 8'h24;
frames[18][19][1] = 8'h24;
frames[18][19][2] = 8'h24;
frames[18][19][3] = 8'h49;
frames[18][19][4] = 8'h48;
frames[18][19][5] = 8'h24;
frames[18][19][6] = 8'h00;
frames[18][19][7] = 8'h6d;
frames[18][19][8] = 8'hff;
frames[18][19][9] = 8'hff;
frames[18][19][10] = 8'hff;
frames[18][19][11] = 8'hff;
frames[18][19][12] = 8'hff;
frames[18][19][13] = 8'hda;
frames[18][19][14] = 8'hb1;
frames[18][19][15] = 8'h68;
frames[18][19][16] = 8'h24;
frames[18][19][17] = 8'h24;
frames[18][19][18] = 8'h24;
frames[18][19][19] = 8'h44;
frames[18][19][20] = 8'h44;
frames[18][19][21] = 8'h44;
frames[18][19][22] = 8'h24;
frames[18][19][23] = 8'h00;
frames[18][19][24] = 8'h00;
frames[18][19][25] = 8'h00;
frames[18][19][26] = 8'h00;
frames[18][19][27] = 8'h20;
frames[18][19][28] = 8'h20;
frames[18][19][29] = 8'h44;
frames[18][19][30] = 8'h48;
frames[18][19][31] = 8'h48;
frames[18][19][32] = 8'h48;
frames[18][19][33] = 8'h24;
frames[18][19][34] = 8'h24;
frames[18][19][35] = 8'h00;
frames[18][19][36] = 8'h00;
frames[18][19][37] = 8'h00;
frames[18][19][38] = 8'h20;
frames[18][19][39] = 8'h20;
frames[18][20][0] = 8'h24;
frames[18][20][1] = 8'h24;
frames[18][20][2] = 8'h00;
frames[18][20][3] = 8'h24;
frames[18][20][4] = 8'h24;
frames[18][20][5] = 8'h49;
frames[18][20][6] = 8'h24;
frames[18][20][7] = 8'h20;
frames[18][20][8] = 8'h8d;
frames[18][20][9] = 8'had;
frames[18][20][10] = 8'had;
frames[18][20][11] = 8'hd1;
frames[18][20][12] = 8'h8d;
frames[18][20][13] = 8'h68;
frames[18][20][14] = 8'h44;
frames[18][20][15] = 8'h20;
frames[18][20][16] = 8'h20;
frames[18][20][17] = 8'h20;
frames[18][20][18] = 8'h20;
frames[18][20][19] = 8'h24;
frames[18][20][20] = 8'h24;
frames[18][20][21] = 8'h00;
frames[18][20][22] = 8'h00;
frames[18][20][23] = 8'h00;
frames[18][20][24] = 8'h00;
frames[18][20][25] = 8'h20;
frames[18][20][26] = 8'h49;
frames[18][20][27] = 8'h49;
frames[18][20][28] = 8'h48;
frames[18][20][29] = 8'h24;
frames[18][20][30] = 8'h04;
frames[18][20][31] = 8'h24;
frames[18][20][32] = 8'h04;
frames[18][20][33] = 8'h28;
frames[18][20][34] = 8'h24;
frames[18][20][35] = 8'h24;
frames[18][20][36] = 8'h24;
frames[18][20][37] = 8'h24;
frames[18][20][38] = 8'h00;
frames[18][20][39] = 8'h00;
frames[18][21][0] = 8'h24;
frames[18][21][1] = 8'h24;
frames[18][21][2] = 8'h04;
frames[18][21][3] = 8'h24;
frames[18][21][4] = 8'h24;
frames[18][21][5] = 8'h24;
frames[18][21][6] = 8'h24;
frames[18][21][7] = 8'h48;
frames[18][21][8] = 8'h44;
frames[18][21][9] = 8'h44;
frames[18][21][10] = 8'h68;
frames[18][21][11] = 8'h68;
frames[18][21][12] = 8'h44;
frames[18][21][13] = 8'h24;
frames[18][21][14] = 8'h00;
frames[18][21][15] = 8'h00;
frames[18][21][16] = 8'h00;
frames[18][21][17] = 8'h00;
frames[18][21][18] = 8'h00;
frames[18][21][19] = 8'h00;
frames[18][21][20] = 8'h00;
frames[18][21][21] = 8'h00;
frames[18][21][22] = 8'h20;
frames[18][21][23] = 8'h20;
frames[18][21][24] = 8'h00;
frames[18][21][25] = 8'h24;
frames[18][21][26] = 8'h6d;
frames[18][21][27] = 8'h71;
frames[18][21][28] = 8'h71;
frames[18][21][29] = 8'h6d;
frames[18][21][30] = 8'h24;
frames[18][21][31] = 8'h6d;
frames[18][21][32] = 8'h28;
frames[18][21][33] = 8'h4d;
frames[18][21][34] = 8'h24;
frames[18][21][35] = 8'h92;
frames[18][21][36] = 8'h92;
frames[18][21][37] = 8'h6d;
frames[18][21][38] = 8'h24;
frames[18][21][39] = 8'h00;
frames[18][22][0] = 8'h20;
frames[18][22][1] = 8'h24;
frames[18][22][2] = 8'h24;
frames[18][22][3] = 8'h24;
frames[18][22][4] = 8'h24;
frames[18][22][5] = 8'h24;
frames[18][22][6] = 8'h24;
frames[18][22][7] = 8'h24;
frames[18][22][8] = 8'h24;
frames[18][22][9] = 8'h44;
frames[18][22][10] = 8'h24;
frames[18][22][11] = 8'h00;
frames[18][22][12] = 8'h00;
frames[18][22][13] = 8'h00;
frames[18][22][14] = 8'h00;
frames[18][22][15] = 8'h00;
frames[18][22][16] = 8'h00;
frames[18][22][17] = 8'h00;
frames[18][22][18] = 8'h00;
frames[18][22][19] = 8'h00;
frames[18][22][20] = 8'h00;
frames[18][22][21] = 8'h24;
frames[18][22][22] = 8'h24;
frames[18][22][23] = 8'h24;
frames[18][22][24] = 8'h24;
frames[18][22][25] = 8'h24;
frames[18][22][26] = 8'h4d;
frames[18][22][27] = 8'h71;
frames[18][22][28] = 8'h71;
frames[18][22][29] = 8'h4d;
frames[18][22][30] = 8'h24;
frames[18][22][31] = 8'h4d;
frames[18][22][32] = 8'h6d;
frames[18][22][33] = 8'h71;
frames[18][22][34] = 8'h49;
frames[18][22][35] = 8'h92;
frames[18][22][36] = 8'h92;
frames[18][22][37] = 8'h92;
frames[18][22][38] = 8'h24;
frames[18][22][39] = 8'h00;
frames[18][23][0] = 8'h20;
frames[18][23][1] = 8'h24;
frames[18][23][2] = 8'h24;
frames[18][23][3] = 8'h24;
frames[18][23][4] = 8'h24;
frames[18][23][5] = 8'h24;
frames[18][23][6] = 8'h24;
frames[18][23][7] = 8'h24;
frames[18][23][8] = 8'h24;
frames[18][23][9] = 8'h24;
frames[18][23][10] = 8'h44;
frames[18][23][11] = 8'h49;
frames[18][23][12] = 8'h48;
frames[18][23][13] = 8'h24;
frames[18][23][14] = 8'h00;
frames[18][23][15] = 8'h00;
frames[18][23][16] = 8'h00;
frames[18][23][17] = 8'h00;
frames[18][23][18] = 8'h00;
frames[18][23][19] = 8'h00;
frames[18][23][20] = 8'h24;
frames[18][23][21] = 8'h24;
frames[18][23][22] = 8'h24;
frames[18][23][23] = 8'h24;
frames[18][23][24] = 8'h24;
frames[18][23][25] = 8'h24;
frames[18][23][26] = 8'h6d;
frames[18][23][27] = 8'h92;
frames[18][23][28] = 8'h71;
frames[18][23][29] = 8'h6d;
frames[18][23][30] = 8'h24;
frames[18][23][31] = 8'h24;
frames[18][23][32] = 8'h28;
frames[18][23][33] = 8'h6d;
frames[18][23][34] = 8'h49;
frames[18][23][35] = 8'h6d;
frames[18][23][36] = 8'h92;
frames[18][23][37] = 8'h92;
frames[18][23][38] = 8'h24;
frames[18][23][39] = 8'h00;
frames[18][24][0] = 8'h00;
frames[18][24][1] = 8'h20;
frames[18][24][2] = 8'h24;
frames[18][24][3] = 8'h24;
frames[18][24][4] = 8'h24;
frames[18][24][5] = 8'h24;
frames[18][24][6] = 8'h24;
frames[18][24][7] = 8'h24;
frames[18][24][8] = 8'h24;
frames[18][24][9] = 8'h24;
frames[18][24][10] = 8'h24;
frames[18][24][11] = 8'h24;
frames[18][24][12] = 8'h49;
frames[18][24][13] = 8'h49;
frames[18][24][14] = 8'h49;
frames[18][24][15] = 8'h24;
frames[18][24][16] = 8'h24;
frames[18][24][17] = 8'h24;
frames[18][24][18] = 8'h24;
frames[18][24][19] = 8'h24;
frames[18][24][20] = 8'h24;
frames[18][24][21] = 8'h24;
frames[18][24][22] = 8'h24;
frames[18][24][23] = 8'h24;
frames[18][24][24] = 8'h24;
frames[18][24][25] = 8'h24;
frames[18][24][26] = 8'h28;
frames[18][24][27] = 8'h24;
frames[18][24][28] = 8'h24;
frames[18][24][29] = 8'h28;
frames[18][24][30] = 8'h24;
frames[18][24][31] = 8'h24;
frames[18][24][32] = 8'h24;
frames[18][24][33] = 8'h24;
frames[18][24][34] = 8'h24;
frames[18][24][35] = 8'h24;
frames[18][24][36] = 8'h24;
frames[18][24][37] = 8'h49;
frames[18][24][38] = 8'h24;
frames[18][24][39] = 8'h24;
frames[18][25][0] = 8'h00;
frames[18][25][1] = 8'h20;
frames[18][25][2] = 8'h24;
frames[18][25][3] = 8'h24;
frames[18][25][4] = 8'h24;
frames[18][25][5] = 8'h24;
frames[18][25][6] = 8'h24;
frames[18][25][7] = 8'h24;
frames[18][25][8] = 8'h24;
frames[18][25][9] = 8'h24;
frames[18][25][10] = 8'h24;
frames[18][25][11] = 8'h24;
frames[18][25][12] = 8'h24;
frames[18][25][13] = 8'h24;
frames[18][25][14] = 8'h49;
frames[18][25][15] = 8'h49;
frames[18][25][16] = 8'h24;
frames[18][25][17] = 8'h24;
frames[18][25][18] = 8'h44;
frames[18][25][19] = 8'h24;
frames[18][25][20] = 8'h24;
frames[18][25][21] = 8'h24;
frames[18][25][22] = 8'h24;
frames[18][25][23] = 8'h24;
frames[18][25][24] = 8'h24;
frames[18][25][25] = 8'h24;
frames[18][25][26] = 8'h6d;
frames[18][25][27] = 8'h6d;
frames[18][25][28] = 8'h6d;
frames[18][25][29] = 8'h71;
frames[18][25][30] = 8'h6d;
frames[18][25][31] = 8'h6d;
frames[18][25][32] = 8'h6d;
frames[18][25][33] = 8'h49;
frames[18][25][34] = 8'h6d;
frames[18][25][35] = 8'h6d;
frames[18][25][36] = 8'h6d;
frames[18][25][37] = 8'h6d;
frames[18][25][38] = 8'h24;
frames[18][25][39] = 8'h24;
frames[18][26][0] = 8'h49;
frames[18][26][1] = 8'h20;
frames[18][26][2] = 8'h00;
frames[18][26][3] = 8'h24;
frames[18][26][4] = 8'h24;
frames[18][26][5] = 8'h24;
frames[18][26][6] = 8'h24;
frames[18][26][7] = 8'h24;
frames[18][26][8] = 8'h24;
frames[18][26][9] = 8'h24;
frames[18][26][10] = 8'h24;
frames[18][26][11] = 8'h24;
frames[18][26][12] = 8'h24;
frames[18][26][13] = 8'h24;
frames[18][26][14] = 8'h24;
frames[18][26][15] = 8'h24;
frames[18][26][16] = 8'h48;
frames[18][26][17] = 8'h49;
frames[18][26][18] = 8'h48;
frames[18][26][19] = 8'h24;
frames[18][26][20] = 8'h24;
frames[18][26][21] = 8'h24;
frames[18][26][22] = 8'h24;
frames[18][26][23] = 8'h24;
frames[18][26][24] = 8'h24;
frames[18][26][25] = 8'h24;
frames[18][26][26] = 8'h49;
frames[18][26][27] = 8'h6d;
frames[18][26][28] = 8'h91;
frames[18][26][29] = 8'h92;
frames[18][26][30] = 8'h92;
frames[18][26][31] = 8'h92;
frames[18][26][32] = 8'h6d;
frames[18][26][33] = 8'h24;
frames[18][26][34] = 8'h4d;
frames[18][26][35] = 8'h92;
frames[18][26][36] = 8'h6d;
frames[18][26][37] = 8'h49;
frames[18][26][38] = 8'h24;
frames[18][26][39] = 8'h04;
frames[18][27][0] = 8'h48;
frames[18][27][1] = 8'h00;
frames[18][27][2] = 8'h00;
frames[18][27][3] = 8'h04;
frames[18][27][4] = 8'h24;
frames[18][27][5] = 8'h24;
frames[18][27][6] = 8'h24;
frames[18][27][7] = 8'h24;
frames[18][27][8] = 8'h24;
frames[18][27][9] = 8'h24;
frames[18][27][10] = 8'h24;
frames[18][27][11] = 8'h24;
frames[18][27][12] = 8'h24;
frames[18][27][13] = 8'h24;
frames[18][27][14] = 8'h24;
frames[18][27][15] = 8'h24;
frames[18][27][16] = 8'h24;
frames[18][27][17] = 8'h24;
frames[18][27][18] = 8'h48;
frames[18][27][19] = 8'h49;
frames[18][27][20] = 8'h48;
frames[18][27][21] = 8'h24;
frames[18][27][22] = 8'h24;
frames[18][27][23] = 8'h24;
frames[18][27][24] = 8'h24;
frames[18][27][25] = 8'h24;
frames[18][27][26] = 8'h49;
frames[18][27][27] = 8'h6d;
frames[18][27][28] = 8'h92;
frames[18][27][29] = 8'h91;
frames[18][27][30] = 8'h92;
frames[18][27][31] = 8'h92;
frames[18][27][32] = 8'h92;
frames[18][27][33] = 8'h49;
frames[18][27][34] = 8'h6d;
frames[18][27][35] = 8'h92;
frames[18][27][36] = 8'h91;
frames[18][27][37] = 8'h6d;
frames[18][27][38] = 8'h24;
frames[18][27][39] = 8'h04;
frames[18][28][0] = 8'h6d;
frames[18][28][1] = 8'h00;
frames[18][28][2] = 8'h00;
frames[18][28][3] = 8'h00;
frames[18][28][4] = 8'h24;
frames[18][28][5] = 8'h24;
frames[18][28][6] = 8'h24;
frames[18][28][7] = 8'h24;
frames[18][28][8] = 8'h24;
frames[18][28][9] = 8'h24;
frames[18][28][10] = 8'h24;
frames[18][28][11] = 8'h24;
frames[18][28][12] = 8'h24;
frames[18][28][13] = 8'h24;
frames[18][28][14] = 8'h24;
frames[18][28][15] = 8'h24;
frames[18][28][16] = 8'h24;
frames[18][28][17] = 8'h24;
frames[18][28][18] = 8'h24;
frames[18][28][19] = 8'h24;
frames[18][28][20] = 8'h48;
frames[18][28][21] = 8'h49;
frames[18][28][22] = 8'h49;
frames[18][28][23] = 8'h44;
frames[18][28][24] = 8'h24;
frames[18][28][25] = 8'h24;
frames[18][28][26] = 8'h24;
frames[18][28][27] = 8'h49;
frames[18][28][28] = 8'h49;
frames[18][28][29] = 8'h49;
frames[18][28][30] = 8'h49;
frames[18][28][31] = 8'h49;
frames[18][28][32] = 8'h49;
frames[18][28][33] = 8'h24;
frames[18][28][34] = 8'h49;
frames[18][28][35] = 8'h49;
frames[18][28][36] = 8'h49;
frames[18][28][37] = 8'h4d;
frames[18][28][38] = 8'h24;
frames[18][28][39] = 8'h00;
frames[18][29][0] = 8'hdb;
frames[18][29][1] = 8'h92;
frames[18][29][2] = 8'h24;
frames[18][29][3] = 8'h24;
frames[18][29][4] = 8'h24;
frames[18][29][5] = 8'h24;
frames[18][29][6] = 8'h24;
frames[18][29][7] = 8'h24;
frames[18][29][8] = 8'h24;
frames[18][29][9] = 8'h24;
frames[18][29][10] = 8'h24;
frames[18][29][11] = 8'h24;
frames[18][29][12] = 8'h24;
frames[18][29][13] = 8'h24;
frames[18][29][14] = 8'h24;
frames[18][29][15] = 8'h24;
frames[18][29][16] = 8'h24;
frames[18][29][17] = 8'h24;
frames[18][29][18] = 8'h24;
frames[18][29][19] = 8'h24;
frames[18][29][20] = 8'h24;
frames[18][29][21] = 8'h24;
frames[18][29][22] = 8'h49;
frames[18][29][23] = 8'h69;
frames[18][29][24] = 8'h49;
frames[18][29][25] = 8'h24;
frames[18][29][26] = 8'h24;
frames[18][29][27] = 8'h00;
frames[18][29][28] = 8'h00;
frames[18][29][29] = 8'h04;
frames[18][29][30] = 8'h04;
frames[18][29][31] = 8'h04;
frames[18][29][32] = 8'h00;
frames[18][29][33] = 8'h24;
frames[18][29][34] = 8'h00;
frames[18][29][35] = 8'h00;
frames[18][29][36] = 8'h00;
frames[18][29][37] = 8'h00;
frames[18][29][38] = 8'h00;
frames[18][29][39] = 8'h04;
frames[19][0][0] = 8'h20;
frames[19][0][1] = 8'h24;
frames[19][0][2] = 8'h91;
frames[19][0][3] = 8'hb6;
frames[19][0][4] = 8'hb6;
frames[19][0][5] = 8'hb6;
frames[19][0][6] = 8'hb6;
frames[19][0][7] = 8'hb6;
frames[19][0][8] = 8'hb1;
frames[19][0][9] = 8'h44;
frames[19][0][10] = 8'h00;
frames[19][0][11] = 8'h00;
frames[19][0][12] = 8'h00;
frames[19][0][13] = 8'h00;
frames[19][0][14] = 8'h00;
frames[19][0][15] = 8'h20;
frames[19][0][16] = 8'h68;
frames[19][0][17] = 8'h91;
frames[19][0][18] = 8'h69;
frames[19][0][19] = 8'h24;
frames[19][0][20] = 8'h00;
frames[19][0][21] = 8'h00;
frames[19][0][22] = 8'h00;
frames[19][0][23] = 8'h24;
frames[19][0][24] = 8'h00;
frames[19][0][25] = 8'h00;
frames[19][0][26] = 8'h00;
frames[19][0][27] = 8'h00;
frames[19][0][28] = 8'h00;
frames[19][0][29] = 8'h00;
frames[19][0][30] = 8'h20;
frames[19][0][31] = 8'h20;
frames[19][0][32] = 8'h20;
frames[19][0][33] = 8'h20;
frames[19][0][34] = 8'h20;
frames[19][0][35] = 8'h20;
frames[19][0][36] = 8'h00;
frames[19][0][37] = 8'h49;
frames[19][0][38] = 8'h24;
frames[19][0][39] = 8'h00;
frames[19][1][0] = 8'h20;
frames[19][1][1] = 8'h24;
frames[19][1][2] = 8'h91;
frames[19][1][3] = 8'hb6;
frames[19][1][4] = 8'hb6;
frames[19][1][5] = 8'hb6;
frames[19][1][6] = 8'hb6;
frames[19][1][7] = 8'hb6;
frames[19][1][8] = 8'hb2;
frames[19][1][9] = 8'h44;
frames[19][1][10] = 8'h00;
frames[19][1][11] = 8'h00;
frames[19][1][12] = 8'h00;
frames[19][1][13] = 8'h00;
frames[19][1][14] = 8'h24;
frames[19][1][15] = 8'h48;
frames[19][1][16] = 8'h6d;
frames[19][1][17] = 8'h48;
frames[19][1][18] = 8'h24;
frames[19][1][19] = 8'h00;
frames[19][1][20] = 8'h00;
frames[19][1][21] = 8'h24;
frames[19][1][22] = 8'h44;
frames[19][1][23] = 8'h20;
frames[19][1][24] = 8'h00;
frames[19][1][25] = 8'h00;
frames[19][1][26] = 8'h00;
frames[19][1][27] = 8'h00;
frames[19][1][28] = 8'h00;
frames[19][1][29] = 8'h00;
frames[19][1][30] = 8'h20;
frames[19][1][31] = 8'h20;
frames[19][1][32] = 8'h24;
frames[19][1][33] = 8'h20;
frames[19][1][34] = 8'h20;
frames[19][1][35] = 8'h20;
frames[19][1][36] = 8'h49;
frames[19][1][37] = 8'hb2;
frames[19][1][38] = 8'hb6;
frames[19][1][39] = 8'h24;
frames[19][2][0] = 8'h20;
frames[19][2][1] = 8'h24;
frames[19][2][2] = 8'h91;
frames[19][2][3] = 8'hb1;
frames[19][2][4] = 8'hb5;
frames[19][2][5] = 8'hb5;
frames[19][2][6] = 8'hb6;
frames[19][2][7] = 8'hb6;
frames[19][2][8] = 8'hb2;
frames[19][2][9] = 8'h68;
frames[19][2][10] = 8'h00;
frames[19][2][11] = 8'h00;
frames[19][2][12] = 8'h00;
frames[19][2][13] = 8'h00;
frames[19][2][14] = 8'h24;
frames[19][2][15] = 8'h6d;
frames[19][2][16] = 8'h48;
frames[19][2][17] = 8'h00;
frames[19][2][18] = 8'h00;
frames[19][2][19] = 8'h00;
frames[19][2][20] = 8'h00;
frames[19][2][21] = 8'h24;
frames[19][2][22] = 8'h48;
frames[19][2][23] = 8'h00;
frames[19][2][24] = 8'h00;
frames[19][2][25] = 8'h00;
frames[19][2][26] = 8'h00;
frames[19][2][27] = 8'h00;
frames[19][2][28] = 8'h00;
frames[19][2][29] = 8'h00;
frames[19][2][30] = 8'h20;
frames[19][2][31] = 8'h24;
frames[19][2][32] = 8'h24;
frames[19][2][33] = 8'h24;
frames[19][2][34] = 8'h24;
frames[19][2][35] = 8'h24;
frames[19][2][36] = 8'h6d;
frames[19][2][37] = 8'h49;
frames[19][2][38] = 8'h4d;
frames[19][2][39] = 8'h4e;
frames[19][3][0] = 8'h20;
frames[19][3][1] = 8'h24;
frames[19][3][2] = 8'h8d;
frames[19][3][3] = 8'hb1;
frames[19][3][4] = 8'hb6;
frames[19][3][5] = 8'hd6;
frames[19][3][6] = 8'hb6;
frames[19][3][7] = 8'hb6;
frames[19][3][8] = 8'hb6;
frames[19][3][9] = 8'h91;
frames[19][3][10] = 8'h24;
frames[19][3][11] = 8'h00;
frames[19][3][12] = 8'h00;
frames[19][3][13] = 8'h00;
frames[19][3][14] = 8'h24;
frames[19][3][15] = 8'h24;
frames[19][3][16] = 8'h04;
frames[19][3][17] = 8'h00;
frames[19][3][18] = 8'h00;
frames[19][3][19] = 8'h00;
frames[19][3][20] = 8'h24;
frames[19][3][21] = 8'h49;
frames[19][3][22] = 8'h24;
frames[19][3][23] = 8'h00;
frames[19][3][24] = 8'h00;
frames[19][3][25] = 8'h00;
frames[19][3][26] = 8'h00;
frames[19][3][27] = 8'h00;
frames[19][3][28] = 8'h00;
frames[19][3][29] = 8'h20;
frames[19][3][30] = 8'h20;
frames[19][3][31] = 8'h24;
frames[19][3][32] = 8'h24;
frames[19][3][33] = 8'h24;
frames[19][3][34] = 8'h24;
frames[19][3][35] = 8'h24;
frames[19][3][36] = 8'h6d;
frames[19][3][37] = 8'h6d;
frames[19][3][38] = 8'h49;
frames[19][3][39] = 8'h6e;
frames[19][4][0] = 8'h00;
frames[19][4][1] = 8'h00;
frames[19][4][2] = 8'h68;
frames[19][4][3] = 8'hb1;
frames[19][4][4] = 8'hd6;
frames[19][4][5] = 8'hb6;
frames[19][4][6] = 8'hb6;
frames[19][4][7] = 8'hb6;
frames[19][4][8] = 8'hb6;
frames[19][4][9] = 8'hb6;
frames[19][4][10] = 8'h6d;
frames[19][4][11] = 8'h00;
frames[19][4][12] = 8'h00;
frames[19][4][13] = 8'h00;
frames[19][4][14] = 8'h00;
frames[19][4][15] = 8'h00;
frames[19][4][16] = 8'h00;
frames[19][4][17] = 8'h24;
frames[19][4][18] = 8'h20;
frames[19][4][19] = 8'h24;
frames[19][4][20] = 8'h6d;
frames[19][4][21] = 8'h24;
frames[19][4][22] = 8'h00;
frames[19][4][23] = 8'h00;
frames[19][4][24] = 8'h00;
frames[19][4][25] = 8'h00;
frames[19][4][26] = 8'h00;
frames[19][4][27] = 8'h00;
frames[19][4][28] = 8'h00;
frames[19][4][29] = 8'h20;
frames[19][4][30] = 8'h24;
frames[19][4][31] = 8'h24;
frames[19][4][32] = 8'h24;
frames[19][4][33] = 8'h24;
frames[19][4][34] = 8'h24;
frames[19][4][35] = 8'h24;
frames[19][4][36] = 8'h92;
frames[19][4][37] = 8'h6d;
frames[19][4][38] = 8'h6e;
frames[19][4][39] = 8'h6e;
frames[19][5][0] = 8'h00;
frames[19][5][1] = 8'h00;
frames[19][5][2] = 8'h48;
frames[19][5][3] = 8'hb2;
frames[19][5][4] = 8'hd6;
frames[19][5][5] = 8'hb6;
frames[19][5][6] = 8'hb6;
frames[19][5][7] = 8'hb6;
frames[19][5][8] = 8'hb6;
frames[19][5][9] = 8'hb5;
frames[19][5][10] = 8'h8d;
frames[19][5][11] = 8'h20;
frames[19][5][12] = 8'h00;
frames[19][5][13] = 8'h00;
frames[19][5][14] = 8'h20;
frames[19][5][15] = 8'h24;
frames[19][5][16] = 8'h20;
frames[19][5][17] = 8'h00;
frames[19][5][18] = 8'h24;
frames[19][5][19] = 8'h6d;
frames[19][5][20] = 8'h49;
frames[19][5][21] = 8'h00;
frames[19][5][22] = 8'h00;
frames[19][5][23] = 8'h00;
frames[19][5][24] = 8'h00;
frames[19][5][25] = 8'h00;
frames[19][5][26] = 8'h00;
frames[19][5][27] = 8'h20;
frames[19][5][28] = 8'h20;
frames[19][5][29] = 8'h24;
frames[19][5][30] = 8'h24;
frames[19][5][31] = 8'h24;
frames[19][5][32] = 8'h24;
frames[19][5][33] = 8'h24;
frames[19][5][34] = 8'h24;
frames[19][5][35] = 8'h24;
frames[19][5][36] = 8'h49;
frames[19][5][37] = 8'h92;
frames[19][5][38] = 8'h92;
frames[19][5][39] = 8'h24;
frames[19][6][0] = 8'h00;
frames[19][6][1] = 8'h00;
frames[19][6][2] = 8'h20;
frames[19][6][3] = 8'h6d;
frames[19][6][4] = 8'hb1;
frames[19][6][5] = 8'hb1;
frames[19][6][6] = 8'hb6;
frames[19][6][7] = 8'hb6;
frames[19][6][8] = 8'hb6;
frames[19][6][9] = 8'hb6;
frames[19][6][10] = 8'hb1;
frames[19][6][11] = 8'h48;
frames[19][6][12] = 8'h00;
frames[19][6][13] = 8'h20;
frames[19][6][14] = 8'h20;
frames[19][6][15] = 8'h20;
frames[19][6][16] = 8'h20;
frames[19][6][17] = 8'h24;
frames[19][6][18] = 8'h8d;
frames[19][6][19] = 8'h6d;
frames[19][6][20] = 8'h24;
frames[19][6][21] = 8'h00;
frames[19][6][22] = 8'h00;
frames[19][6][23] = 8'h00;
frames[19][6][24] = 8'h00;
frames[19][6][25] = 8'h00;
frames[19][6][26] = 8'h00;
frames[19][6][27] = 8'h24;
frames[19][6][28] = 8'h24;
frames[19][6][29] = 8'h24;
frames[19][6][30] = 8'h24;
frames[19][6][31] = 8'h24;
frames[19][6][32] = 8'h24;
frames[19][6][33] = 8'h24;
frames[19][6][34] = 8'h24;
frames[19][6][35] = 8'h24;
frames[19][6][36] = 8'h24;
frames[19][6][37] = 8'h24;
frames[19][6][38] = 8'h24;
frames[19][6][39] = 8'h24;
frames[19][7][0] = 8'h24;
frames[19][7][1] = 8'h24;
frames[19][7][2] = 8'h48;
frames[19][7][3] = 8'h8d;
frames[19][7][4] = 8'h91;
frames[19][7][5] = 8'hb1;
frames[19][7][6] = 8'hb6;
frames[19][7][7] = 8'hb6;
frames[19][7][8] = 8'hb6;
frames[19][7][9] = 8'hb6;
frames[19][7][10] = 8'hb1;
frames[19][7][11] = 8'h8d;
frames[19][7][12] = 8'h20;
frames[19][7][13] = 8'h00;
frames[19][7][14] = 8'h00;
frames[19][7][15] = 8'h00;
frames[19][7][16] = 8'h20;
frames[19][7][17] = 8'h49;
frames[19][7][18] = 8'h8d;
frames[19][7][19] = 8'h44;
frames[19][7][20] = 8'h00;
frames[19][7][21] = 8'h00;
frames[19][7][22] = 8'h00;
frames[19][7][23] = 8'h00;
frames[19][7][24] = 8'h00;
frames[19][7][25] = 8'h00;
frames[19][7][26] = 8'h20;
frames[19][7][27] = 8'h24;
frames[19][7][28] = 8'h24;
frames[19][7][29] = 8'h24;
frames[19][7][30] = 8'h24;
frames[19][7][31] = 8'h24;
frames[19][7][32] = 8'h24;
frames[19][7][33] = 8'h24;
frames[19][7][34] = 8'h24;
frames[19][7][35] = 8'h24;
frames[19][7][36] = 8'h24;
frames[19][7][37] = 8'h24;
frames[19][7][38] = 8'h24;
frames[19][7][39] = 8'h24;
frames[19][8][0] = 8'hd6;
frames[19][8][1] = 8'hda;
frames[19][8][2] = 8'hda;
frames[19][8][3] = 8'hda;
frames[19][8][4] = 8'h8d;
frames[19][8][5] = 8'h8d;
frames[19][8][6] = 8'hb5;
frames[19][8][7] = 8'hb5;
frames[19][8][8] = 8'hb6;
frames[19][8][9] = 8'hb6;
frames[19][8][10] = 8'hb6;
frames[19][8][11] = 8'hb5;
frames[19][8][12] = 8'h48;
frames[19][8][13] = 8'h00;
frames[19][8][14] = 8'h00;
frames[19][8][15] = 8'h00;
frames[19][8][16] = 8'h00;
frames[19][8][17] = 8'h24;
frames[19][8][18] = 8'h24;
frames[19][8][19] = 8'h24;
frames[19][8][20] = 8'h00;
frames[19][8][21] = 8'h00;
frames[19][8][22] = 8'h00;
frames[19][8][23] = 8'h00;
frames[19][8][24] = 8'h00;
frames[19][8][25] = 8'h00;
frames[19][8][26] = 8'h20;
frames[19][8][27] = 8'h24;
frames[19][8][28] = 8'h24;
frames[19][8][29] = 8'h24;
frames[19][8][30] = 8'h24;
frames[19][8][31] = 8'h24;
frames[19][8][32] = 8'h24;
frames[19][8][33] = 8'h24;
frames[19][8][34] = 8'h24;
frames[19][8][35] = 8'h24;
frames[19][8][36] = 8'h24;
frames[19][8][37] = 8'h24;
frames[19][8][38] = 8'h24;
frames[19][8][39] = 8'h24;
frames[19][9][0] = 8'hfa;
frames[19][9][1] = 8'hda;
frames[19][9][2] = 8'hda;
frames[19][9][3] = 8'hfa;
frames[19][9][4] = 8'hb1;
frames[19][9][5] = 8'h8d;
frames[19][9][6] = 8'hb1;
frames[19][9][7] = 8'hb6;
frames[19][9][8] = 8'hb6;
frames[19][9][9] = 8'hb6;
frames[19][9][10] = 8'hb6;
frames[19][9][11] = 8'hb6;
frames[19][9][12] = 8'h6d;
frames[19][9][13] = 8'h20;
frames[19][9][14] = 8'h20;
frames[19][9][15] = 8'h20;
frames[19][9][16] = 8'h20;
frames[19][9][17] = 8'h20;
frames[19][9][18] = 8'h00;
frames[19][9][19] = 8'h00;
frames[19][9][20] = 8'h00;
frames[19][9][21] = 8'h00;
frames[19][9][22] = 8'h00;
frames[19][9][23] = 8'h00;
frames[19][9][24] = 8'h00;
frames[19][9][25] = 8'h20;
frames[19][9][26] = 8'h24;
frames[19][9][27] = 8'h24;
frames[19][9][28] = 8'h24;
frames[19][9][29] = 8'h24;
frames[19][9][30] = 8'h24;
frames[19][9][31] = 8'h24;
frames[19][9][32] = 8'h24;
frames[19][9][33] = 8'h24;
frames[19][9][34] = 8'h24;
frames[19][9][35] = 8'h24;
frames[19][9][36] = 8'h24;
frames[19][9][37] = 8'h24;
frames[19][9][38] = 8'h24;
frames[19][9][39] = 8'h24;
frames[19][10][0] = 8'hda;
frames[19][10][1] = 8'hda;
frames[19][10][2] = 8'hda;
frames[19][10][3] = 8'hda;
frames[19][10][4] = 8'hb6;
frames[19][10][5] = 8'h6d;
frames[19][10][6] = 8'h91;
frames[19][10][7] = 8'hd6;
frames[19][10][8] = 8'hd6;
frames[19][10][9] = 8'hb6;
frames[19][10][10] = 8'hb6;
frames[19][10][11] = 8'hb6;
frames[19][10][12] = 8'hb6;
frames[19][10][13] = 8'h48;
frames[19][10][14] = 8'h24;
frames[19][10][15] = 8'h20;
frames[19][10][16] = 8'h00;
frames[19][10][17] = 8'h00;
frames[19][10][18] = 8'h00;
frames[19][10][19] = 8'h00;
frames[19][10][20] = 8'h00;
frames[19][10][21] = 8'h00;
frames[19][10][22] = 8'h00;
frames[19][10][23] = 8'h00;
frames[19][10][24] = 8'h20;
frames[19][10][25] = 8'h20;
frames[19][10][26] = 8'h24;
frames[19][10][27] = 8'h20;
frames[19][10][28] = 8'h24;
frames[19][10][29] = 8'h24;
frames[19][10][30] = 8'h24;
frames[19][10][31] = 8'h24;
frames[19][10][32] = 8'h24;
frames[19][10][33] = 8'h20;
frames[19][10][34] = 8'h20;
frames[19][10][35] = 8'h20;
frames[19][10][36] = 8'h20;
frames[19][10][37] = 8'h20;
frames[19][10][38] = 8'h20;
frames[19][10][39] = 8'h00;
frames[19][11][0] = 8'hda;
frames[19][11][1] = 8'hda;
frames[19][11][2] = 8'hda;
frames[19][11][3] = 8'hfa;
frames[19][11][4] = 8'hda;
frames[19][11][5] = 8'h8d;
frames[19][11][6] = 8'h8d;
frames[19][11][7] = 8'hb6;
frames[19][11][8] = 8'hd6;
frames[19][11][9] = 8'hd6;
frames[19][11][10] = 8'hd6;
frames[19][11][11] = 8'hb6;
frames[19][11][12] = 8'hd6;
frames[19][11][13] = 8'h8d;
frames[19][11][14] = 8'h24;
frames[19][11][15] = 8'h20;
frames[19][11][16] = 8'h20;
frames[19][11][17] = 8'h20;
frames[19][11][18] = 8'h24;
frames[19][11][19] = 8'h20;
frames[19][11][20] = 8'h00;
frames[19][11][21] = 8'h00;
frames[19][11][22] = 8'h00;
frames[19][11][23] = 8'h00;
frames[19][11][24] = 8'h00;
frames[19][11][25] = 8'h00;
frames[19][11][26] = 8'h00;
frames[19][11][27] = 8'h00;
frames[19][11][28] = 8'h20;
frames[19][11][29] = 8'h24;
frames[19][11][30] = 8'h24;
frames[19][11][31] = 8'h24;
frames[19][11][32] = 8'h24;
frames[19][11][33] = 8'h20;
frames[19][11][34] = 8'h00;
frames[19][11][35] = 8'h20;
frames[19][11][36] = 8'h00;
frames[19][11][37] = 8'h20;
frames[19][11][38] = 8'h20;
frames[19][11][39] = 8'h24;
frames[19][12][0] = 8'hfa;
frames[19][12][1] = 8'hfa;
frames[19][12][2] = 8'hfa;
frames[19][12][3] = 8'hfa;
frames[19][12][4] = 8'hfb;
frames[19][12][5] = 8'hd6;
frames[19][12][6] = 8'h8d;
frames[19][12][7] = 8'h91;
frames[19][12][8] = 8'hb6;
frames[19][12][9] = 8'hb6;
frames[19][12][10] = 8'hb5;
frames[19][12][11] = 8'hb1;
frames[19][12][12] = 8'hb6;
frames[19][12][13] = 8'hb1;
frames[19][12][14] = 8'h48;
frames[19][12][15] = 8'h00;
frames[19][12][16] = 8'h00;
frames[19][12][17] = 8'h20;
frames[19][12][18] = 8'h20;
frames[19][12][19] = 8'h00;
frames[19][12][20] = 8'h00;
frames[19][12][21] = 8'h00;
frames[19][12][22] = 8'h20;
frames[19][12][23] = 8'h24;
frames[19][12][24] = 8'h24;
frames[19][12][25] = 8'h20;
frames[19][12][26] = 8'h00;
frames[19][12][27] = 8'h00;
frames[19][12][28] = 8'h00;
frames[19][12][29] = 8'h00;
frames[19][12][30] = 8'h00;
frames[19][12][31] = 8'h00;
frames[19][12][32] = 8'h00;
frames[19][12][33] = 8'h00;
frames[19][12][34] = 8'h00;
frames[19][12][35] = 8'h00;
frames[19][12][36] = 8'h00;
frames[19][12][37] = 8'h00;
frames[19][12][38] = 8'h24;
frames[19][12][39] = 8'h20;
frames[19][13][0] = 8'hfa;
frames[19][13][1] = 8'hfa;
frames[19][13][2] = 8'hfb;
frames[19][13][3] = 8'hfa;
frames[19][13][4] = 8'hd6;
frames[19][13][5] = 8'hb1;
frames[19][13][6] = 8'h8d;
frames[19][13][7] = 8'h8d;
frames[19][13][8] = 8'hb1;
frames[19][13][9] = 8'hb1;
frames[19][13][10] = 8'hb6;
frames[19][13][11] = 8'hb6;
frames[19][13][12] = 8'hd6;
frames[19][13][13] = 8'hb6;
frames[19][13][14] = 8'h91;
frames[19][13][15] = 8'h24;
frames[19][13][16] = 8'h00;
frames[19][13][17] = 8'h00;
frames[19][13][18] = 8'h00;
frames[19][13][19] = 8'h00;
frames[19][13][20] = 8'h00;
frames[19][13][21] = 8'h24;
frames[19][13][22] = 8'h24;
frames[19][13][23] = 8'h24;
frames[19][13][24] = 8'h24;
frames[19][13][25] = 8'h20;
frames[19][13][26] = 8'h00;
frames[19][13][27] = 8'h00;
frames[19][13][28] = 8'h00;
frames[19][13][29] = 8'h00;
frames[19][13][30] = 8'h00;
frames[19][13][31] = 8'h00;
frames[19][13][32] = 8'h00;
frames[19][13][33] = 8'h00;
frames[19][13][34] = 8'h00;
frames[19][13][35] = 8'h00;
frames[19][13][36] = 8'h24;
frames[19][13][37] = 8'h24;
frames[19][13][38] = 8'h24;
frames[19][13][39] = 8'h00;
frames[19][14][0] = 8'hd6;
frames[19][14][1] = 8'hb1;
frames[19][14][2] = 8'h8d;
frames[19][14][3] = 8'h68;
frames[19][14][4] = 8'h44;
frames[19][14][5] = 8'h44;
frames[19][14][6] = 8'h44;
frames[19][14][7] = 8'h48;
frames[19][14][8] = 8'h68;
frames[19][14][9] = 8'hb1;
frames[19][14][10] = 8'hb5;
frames[19][14][11] = 8'hd6;
frames[19][14][12] = 8'hd6;
frames[19][14][13] = 8'hd6;
frames[19][14][14] = 8'hd6;
frames[19][14][15] = 8'hb2;
frames[19][14][16] = 8'h6d;
frames[19][14][17] = 8'h69;
frames[19][14][18] = 8'h48;
frames[19][14][19] = 8'h49;
frames[19][14][20] = 8'h69;
frames[19][14][21] = 8'h44;
frames[19][14][22] = 8'h20;
frames[19][14][23] = 8'h00;
frames[19][14][24] = 8'h00;
frames[19][14][25] = 8'h00;
frames[19][14][26] = 8'h00;
frames[19][14][27] = 8'h00;
frames[19][14][28] = 8'h00;
frames[19][14][29] = 8'h00;
frames[19][14][30] = 8'h00;
frames[19][14][31] = 8'h00;
frames[19][14][32] = 8'h00;
frames[19][14][33] = 8'h00;
frames[19][14][34] = 8'h24;
frames[19][14][35] = 8'h24;
frames[19][14][36] = 8'h24;
frames[19][14][37] = 8'h00;
frames[19][14][38] = 8'h00;
frames[19][14][39] = 8'h00;
frames[19][15][0] = 8'h44;
frames[19][15][1] = 8'h24;
frames[19][15][2] = 8'h20;
frames[19][15][3] = 8'h00;
frames[19][15][4] = 8'h00;
frames[19][15][5] = 8'h00;
frames[19][15][6] = 8'h00;
frames[19][15][7] = 8'h00;
frames[19][15][8] = 8'h24;
frames[19][15][9] = 8'h69;
frames[19][15][10] = 8'hb1;
frames[19][15][11] = 8'hb6;
frames[19][15][12] = 8'hd6;
frames[19][15][13] = 8'hd6;
frames[19][15][14] = 8'hd6;
frames[19][15][15] = 8'hd6;
frames[19][15][16] = 8'hd6;
frames[19][15][17] = 8'hb6;
frames[19][15][18] = 8'h91;
frames[19][15][19] = 8'h8d;
frames[19][15][20] = 8'h49;
frames[19][15][21] = 8'h24;
frames[19][15][22] = 8'h00;
frames[19][15][23] = 8'h00;
frames[19][15][24] = 8'h00;
frames[19][15][25] = 8'h00;
frames[19][15][26] = 8'h00;
frames[19][15][27] = 8'h00;
frames[19][15][28] = 8'h00;
frames[19][15][29] = 8'h00;
frames[19][15][30] = 8'h00;
frames[19][15][31] = 8'h00;
frames[19][15][32] = 8'h00;
frames[19][15][33] = 8'h24;
frames[19][15][34] = 8'h24;
frames[19][15][35] = 8'h24;
frames[19][15][36] = 8'h00;
frames[19][15][37] = 8'h00;
frames[19][15][38] = 8'h00;
frames[19][15][39] = 8'h00;
frames[19][16][0] = 8'h20;
frames[19][16][1] = 8'h00;
frames[19][16][2] = 8'h00;
frames[19][16][3] = 8'h00;
frames[19][16][4] = 8'h00;
frames[19][16][5] = 8'h00;
frames[19][16][6] = 8'h00;
frames[19][16][7] = 8'h00;
frames[19][16][8] = 8'h20;
frames[19][16][9] = 8'h24;
frames[19][16][10] = 8'h48;
frames[19][16][11] = 8'h6d;
frames[19][16][12] = 8'h91;
frames[19][16][13] = 8'hb1;
frames[19][16][14] = 8'hd6;
frames[19][16][15] = 8'hd6;
frames[19][16][16] = 8'hb6;
frames[19][16][17] = 8'h91;
frames[19][16][18] = 8'h68;
frames[19][16][19] = 8'h24;
frames[19][16][20] = 8'h20;
frames[19][16][21] = 8'h00;
frames[19][16][22] = 8'h00;
frames[19][16][23] = 8'h00;
frames[19][16][24] = 8'h00;
frames[19][16][25] = 8'h00;
frames[19][16][26] = 8'h00;
frames[19][16][27] = 8'h00;
frames[19][16][28] = 8'h00;
frames[19][16][29] = 8'h00;
frames[19][16][30] = 8'h00;
frames[19][16][31] = 8'h20;
frames[19][16][32] = 8'h24;
frames[19][16][33] = 8'h24;
frames[19][16][34] = 8'h00;
frames[19][16][35] = 8'h00;
frames[19][16][36] = 8'h00;
frames[19][16][37] = 8'h00;
frames[19][16][38] = 8'h00;
frames[19][16][39] = 8'h00;
frames[19][17][0] = 8'h20;
frames[19][17][1] = 8'h00;
frames[19][17][2] = 8'h00;
frames[19][17][3] = 8'h20;
frames[19][17][4] = 8'h20;
frames[19][17][5] = 8'h20;
frames[19][17][6] = 8'h20;
frames[19][17][7] = 8'h20;
frames[19][17][8] = 8'h00;
frames[19][17][9] = 8'h00;
frames[19][17][10] = 8'h00;
frames[19][17][11] = 8'h24;
frames[19][17][12] = 8'h24;
frames[19][17][13] = 8'h48;
frames[19][17][14] = 8'h69;
frames[19][17][15] = 8'h48;
frames[19][17][16] = 8'h48;
frames[19][17][17] = 8'h24;
frames[19][17][18] = 8'h00;
frames[19][17][19] = 8'h00;
frames[19][17][20] = 8'h00;
frames[19][17][21] = 8'h00;
frames[19][17][22] = 8'h00;
frames[19][17][23] = 8'h00;
frames[19][17][24] = 8'h00;
frames[19][17][25] = 8'h00;
frames[19][17][26] = 8'h00;
frames[19][17][27] = 8'h00;
frames[19][17][28] = 8'h00;
frames[19][17][29] = 8'h00;
frames[19][17][30] = 8'h24;
frames[19][17][31] = 8'h24;
frames[19][17][32] = 8'h20;
frames[19][17][33] = 8'h20;
frames[19][17][34] = 8'h00;
frames[19][17][35] = 8'h00;
frames[19][17][36] = 8'h00;
frames[19][17][37] = 8'h00;
frames[19][17][38] = 8'h00;
frames[19][17][39] = 8'h00;
frames[19][18][0] = 8'h24;
frames[19][18][1] = 8'h00;
frames[19][18][2] = 8'h20;
frames[19][18][3] = 8'h20;
frames[19][18][4] = 8'h24;
frames[19][18][5] = 8'h24;
frames[19][18][6] = 8'h00;
frames[19][18][7] = 8'h00;
frames[19][18][8] = 8'h00;
frames[19][18][9] = 8'h00;
frames[19][18][10] = 8'h00;
frames[19][18][11] = 8'h00;
frames[19][18][12] = 8'h00;
frames[19][18][13] = 8'h20;
frames[19][18][14] = 8'h20;
frames[19][18][15] = 8'h00;
frames[19][18][16] = 8'h00;
frames[19][18][17] = 8'h00;
frames[19][18][18] = 8'h00;
frames[19][18][19] = 8'h00;
frames[19][18][20] = 8'h00;
frames[19][18][21] = 8'h00;
frames[19][18][22] = 8'h00;
frames[19][18][23] = 8'h00;
frames[19][18][24] = 8'h00;
frames[19][18][25] = 8'h00;
frames[19][18][26] = 8'h20;
frames[19][18][27] = 8'h00;
frames[19][18][28] = 8'h20;
frames[19][18][29] = 8'h24;
frames[19][18][30] = 8'h24;
frames[19][18][31] = 8'h20;
frames[19][18][32] = 8'h00;
frames[19][18][33] = 8'h00;
frames[19][18][34] = 8'h00;
frames[19][18][35] = 8'h00;
frames[19][18][36] = 8'h00;
frames[19][18][37] = 8'h00;
frames[19][18][38] = 8'h00;
frames[19][18][39] = 8'h00;
frames[19][19][0] = 8'h24;
frames[19][19][1] = 8'h20;
frames[19][19][2] = 8'h20;
frames[19][19][3] = 8'h20;
frames[19][19][4] = 8'h24;
frames[19][19][5] = 8'h24;
frames[19][19][6] = 8'h00;
frames[19][19][7] = 8'h00;
frames[19][19][8] = 8'h00;
frames[19][19][9] = 8'h00;
frames[19][19][10] = 8'h00;
frames[19][19][11] = 8'h00;
frames[19][19][12] = 8'h20;
frames[19][19][13] = 8'h20;
frames[19][19][14] = 8'h20;
frames[19][19][15] = 8'h00;
frames[19][19][16] = 8'h00;
frames[19][19][17] = 8'h00;
frames[19][19][18] = 8'h00;
frames[19][19][19] = 8'h00;
frames[19][19][20] = 8'h24;
frames[19][19][21] = 8'h20;
frames[19][19][22] = 8'h24;
frames[19][19][23] = 8'h24;
frames[19][19][24] = 8'h24;
frames[19][19][25] = 8'h24;
frames[19][19][26] = 8'h20;
frames[19][19][27] = 8'h24;
frames[19][19][28] = 8'h24;
frames[19][19][29] = 8'h24;
frames[19][19][30] = 8'h24;
frames[19][19][31] = 8'h00;
frames[19][19][32] = 8'h00;
frames[19][19][33] = 8'h00;
frames[19][19][34] = 8'h00;
frames[19][19][35] = 8'h00;
frames[19][19][36] = 8'h00;
frames[19][19][37] = 8'h00;
frames[19][19][38] = 8'h00;
frames[19][19][39] = 8'h00;
frames[19][20][0] = 8'h44;
frames[19][20][1] = 8'h24;
frames[19][20][2] = 8'h20;
frames[19][20][3] = 8'h20;
frames[19][20][4] = 8'h20;
frames[19][20][5] = 8'h20;
frames[19][20][6] = 8'h00;
frames[19][20][7] = 8'h00;
frames[19][20][8] = 8'h00;
frames[19][20][9] = 8'h00;
frames[19][20][10] = 8'h00;
frames[19][20][11] = 8'h00;
frames[19][20][12] = 8'h20;
frames[19][20][13] = 8'h20;
frames[19][20][14] = 8'h20;
frames[19][20][15] = 8'h20;
frames[19][20][16] = 8'h20;
frames[19][20][17] = 8'h20;
frames[19][20][18] = 8'h24;
frames[19][20][19] = 8'h24;
frames[19][20][20] = 8'h24;
frames[19][20][21] = 8'h24;
frames[19][20][22] = 8'h24;
frames[19][20][23] = 8'h24;
frames[19][20][24] = 8'h24;
frames[19][20][25] = 8'h24;
frames[19][20][26] = 8'h49;
frames[19][20][27] = 8'h49;
frames[19][20][28] = 8'h49;
frames[19][20][29] = 8'h24;
frames[19][20][30] = 8'h24;
frames[19][20][31] = 8'h44;
frames[19][20][32] = 8'h24;
frames[19][20][33] = 8'h44;
frames[19][20][34] = 8'h24;
frames[19][20][35] = 8'h24;
frames[19][20][36] = 8'h44;
frames[19][20][37] = 8'h44;
frames[19][20][38] = 8'h24;
frames[19][20][39] = 8'h00;
frames[19][21][0] = 8'h44;
frames[19][21][1] = 8'h24;
frames[19][21][2] = 8'h20;
frames[19][21][3] = 8'h00;
frames[19][21][4] = 8'h00;
frames[19][21][5] = 8'h00;
frames[19][21][6] = 8'h00;
frames[19][21][7] = 8'h00;
frames[19][21][8] = 8'h00;
frames[19][21][9] = 8'h00;
frames[19][21][10] = 8'h00;
frames[19][21][11] = 8'h00;
frames[19][21][12] = 8'h00;
frames[19][21][13] = 8'h20;
frames[19][21][14] = 8'h20;
frames[19][21][15] = 8'h20;
frames[19][21][16] = 8'h20;
frames[19][21][17] = 8'h20;
frames[19][21][18] = 8'h20;
frames[19][21][19] = 8'h20;
frames[19][21][20] = 8'h20;
frames[19][21][21] = 8'h24;
frames[19][21][22] = 8'h24;
frames[19][21][23] = 8'h24;
frames[19][21][24] = 8'h24;
frames[19][21][25] = 8'h24;
frames[19][21][26] = 8'h69;
frames[19][21][27] = 8'h8d;
frames[19][21][28] = 8'h92;
frames[19][21][29] = 8'h69;
frames[19][21][30] = 8'h24;
frames[19][21][31] = 8'h6d;
frames[19][21][32] = 8'h44;
frames[19][21][33] = 8'h69;
frames[19][21][34] = 8'h24;
frames[19][21][35] = 8'hb2;
frames[19][21][36] = 8'h92;
frames[19][21][37] = 8'h8e;
frames[19][21][38] = 8'h24;
frames[19][21][39] = 8'h00;
frames[19][22][0] = 8'h44;
frames[19][22][1] = 8'h44;
frames[19][22][2] = 8'h20;
frames[19][22][3] = 8'h00;
frames[19][22][4] = 8'h00;
frames[19][22][5] = 8'h00;
frames[19][22][6] = 8'h00;
frames[19][22][7] = 8'h00;
frames[19][22][8] = 8'h00;
frames[19][22][9] = 8'h00;
frames[19][22][10] = 8'h00;
frames[19][22][11] = 8'h00;
frames[19][22][12] = 8'h20;
frames[19][22][13] = 8'h20;
frames[19][22][14] = 8'h20;
frames[19][22][15] = 8'h00;
frames[19][22][16] = 8'h00;
frames[19][22][17] = 8'h20;
frames[19][22][18] = 8'h00;
frames[19][22][19] = 8'h20;
frames[19][22][20] = 8'h20;
frames[19][22][21] = 8'h24;
frames[19][22][22] = 8'h24;
frames[19][22][23] = 8'h24;
frames[19][22][24] = 8'h24;
frames[19][22][25] = 8'h24;
frames[19][22][26] = 8'h69;
frames[19][22][27] = 8'h92;
frames[19][22][28] = 8'h8d;
frames[19][22][29] = 8'h49;
frames[19][22][30] = 8'h24;
frames[19][22][31] = 8'h69;
frames[19][22][32] = 8'h6d;
frames[19][22][33] = 8'h8d;
frames[19][22][34] = 8'h49;
frames[19][22][35] = 8'h92;
frames[19][22][36] = 8'h92;
frames[19][22][37] = 8'h92;
frames[19][22][38] = 8'h24;
frames[19][22][39] = 8'h00;
frames[19][23][0] = 8'h44;
frames[19][23][1] = 8'h48;
frames[19][23][2] = 8'h24;
frames[19][23][3] = 8'h00;
frames[19][23][4] = 8'h00;
frames[19][23][5] = 8'h00;
frames[19][23][6] = 8'h00;
frames[19][23][7] = 8'h00;
frames[19][23][8] = 8'h00;
frames[19][23][9] = 8'h20;
frames[19][23][10] = 8'h24;
frames[19][23][11] = 8'h24;
frames[19][23][12] = 8'h24;
frames[19][23][13] = 8'h24;
frames[19][23][14] = 8'h20;
frames[19][23][15] = 8'h20;
frames[19][23][16] = 8'h20;
frames[19][23][17] = 8'h20;
frames[19][23][18] = 8'h20;
frames[19][23][19] = 8'h20;
frames[19][23][20] = 8'h24;
frames[19][23][21] = 8'h24;
frames[19][23][22] = 8'h24;
frames[19][23][23] = 8'h24;
frames[19][23][24] = 8'h24;
frames[19][23][25] = 8'h24;
frames[19][23][26] = 8'h6d;
frames[19][23][27] = 8'h92;
frames[19][23][28] = 8'h91;
frames[19][23][29] = 8'h6d;
frames[19][23][30] = 8'h49;
frames[19][23][31] = 8'h24;
frames[19][23][32] = 8'h44;
frames[19][23][33] = 8'h6d;
frames[19][23][34] = 8'h49;
frames[19][23][35] = 8'h49;
frames[19][23][36] = 8'h6d;
frames[19][23][37] = 8'h92;
frames[19][23][38] = 8'h24;
frames[19][23][39] = 8'h00;
frames[19][24][0] = 8'h44;
frames[19][24][1] = 8'h44;
frames[19][24][2] = 8'h44;
frames[19][24][3] = 8'h24;
frames[19][24][4] = 8'h24;
frames[19][24][5] = 8'h24;
frames[19][24][6] = 8'h24;
frames[19][24][7] = 8'h24;
frames[19][24][8] = 8'h24;
frames[19][24][9] = 8'h24;
frames[19][24][10] = 8'h24;
frames[19][24][11] = 8'h24;
frames[19][24][12] = 8'h24;
frames[19][24][13] = 8'h24;
frames[19][24][14] = 8'h20;
frames[19][24][15] = 8'h24;
frames[19][24][16] = 8'h24;
frames[19][24][17] = 8'h24;
frames[19][24][18] = 8'h24;
frames[19][24][19] = 8'h24;
frames[19][24][20] = 8'h24;
frames[19][24][21] = 8'h24;
frames[19][24][22] = 8'h24;
frames[19][24][23] = 8'h20;
frames[19][24][24] = 8'h20;
frames[19][24][25] = 8'h20;
frames[19][24][26] = 8'h24;
frames[19][24][27] = 8'h24;
frames[19][24][28] = 8'h24;
frames[19][24][29] = 8'h48;
frames[19][24][30] = 8'h24;
frames[19][24][31] = 8'h24;
frames[19][24][32] = 8'h24;
frames[19][24][33] = 8'h24;
frames[19][24][34] = 8'h24;
frames[19][24][35] = 8'h24;
frames[19][24][36] = 8'h24;
frames[19][24][37] = 8'h24;
frames[19][24][38] = 8'h24;
frames[19][24][39] = 8'h00;
frames[19][25][0] = 8'h24;
frames[19][25][1] = 8'h24;
frames[19][25][2] = 8'h24;
frames[19][25][3] = 8'h44;
frames[19][25][4] = 8'h48;
frames[19][25][5] = 8'h48;
frames[19][25][6] = 8'h48;
frames[19][25][7] = 8'h48;
frames[19][25][8] = 8'h48;
frames[19][25][9] = 8'h44;
frames[19][25][10] = 8'h44;
frames[19][25][11] = 8'h44;
frames[19][25][12] = 8'h24;
frames[19][25][13] = 8'h24;
frames[19][25][14] = 8'h24;
frames[19][25][15] = 8'h24;
frames[19][25][16] = 8'h24;
frames[19][25][17] = 8'h24;
frames[19][25][18] = 8'h24;
frames[19][25][19] = 8'h24;
frames[19][25][20] = 8'h24;
frames[19][25][21] = 8'h24;
frames[19][25][22] = 8'h20;
frames[19][25][23] = 8'h00;
frames[19][25][24] = 8'h00;
frames[19][25][25] = 8'h20;
frames[19][25][26] = 8'h69;
frames[19][25][27] = 8'h6d;
frames[19][25][28] = 8'h6d;
frames[19][25][29] = 8'h8d;
frames[19][25][30] = 8'h6d;
frames[19][25][31] = 8'h91;
frames[19][25][32] = 8'h6d;
frames[19][25][33] = 8'h49;
frames[19][25][34] = 8'h6d;
frames[19][25][35] = 8'h6d;
frames[19][25][36] = 8'h6d;
frames[19][25][37] = 8'h6d;
frames[19][25][38] = 8'h24;
frames[19][25][39] = 8'h00;
frames[19][26][0] = 8'h24;
frames[19][26][1] = 8'h24;
frames[19][26][2] = 8'h24;
frames[19][26][3] = 8'h24;
frames[19][26][4] = 8'h24;
frames[19][26][5] = 8'h24;
frames[19][26][6] = 8'h24;
frames[19][26][7] = 8'h24;
frames[19][26][8] = 8'h24;
frames[19][26][9] = 8'h24;
frames[19][26][10] = 8'h44;
frames[19][26][11] = 8'h44;
frames[19][26][12] = 8'h48;
frames[19][26][13] = 8'h48;
frames[19][26][14] = 8'h48;
frames[19][26][15] = 8'h48;
frames[19][26][16] = 8'h44;
frames[19][26][17] = 8'h24;
frames[19][26][18] = 8'h24;
frames[19][26][19] = 8'h24;
frames[19][26][20] = 8'h20;
frames[19][26][21] = 8'h20;
frames[19][26][22] = 8'h00;
frames[19][26][23] = 8'h00;
frames[19][26][24] = 8'h00;
frames[19][26][25] = 8'h00;
frames[19][26][26] = 8'h44;
frames[19][26][27] = 8'h6d;
frames[19][26][28] = 8'h92;
frames[19][26][29] = 8'h92;
frames[19][26][30] = 8'h92;
frames[19][26][31] = 8'h92;
frames[19][26][32] = 8'h6d;
frames[19][26][33] = 8'h24;
frames[19][26][34] = 8'h6d;
frames[19][26][35] = 8'h92;
frames[19][26][36] = 8'h6d;
frames[19][26][37] = 8'h49;
frames[19][26][38] = 8'h24;
frames[19][26][39] = 8'h00;
frames[19][27][0] = 8'h24;
frames[19][27][1] = 8'h24;
frames[19][27][2] = 8'h24;
frames[19][27][3] = 8'h24;
frames[19][27][4] = 8'h24;
frames[19][27][5] = 8'h24;
frames[19][27][6] = 8'h24;
frames[19][27][7] = 8'h24;
frames[19][27][8] = 8'h24;
frames[19][27][9] = 8'h24;
frames[19][27][10] = 8'h24;
frames[19][27][11] = 8'h24;
frames[19][27][12] = 8'h24;
frames[19][27][13] = 8'h24;
frames[19][27][14] = 8'h24;
frames[19][27][15] = 8'h24;
frames[19][27][16] = 8'h24;
frames[19][27][17] = 8'h24;
frames[19][27][18] = 8'h24;
frames[19][27][19] = 8'h20;
frames[19][27][20] = 8'h00;
frames[19][27][21] = 8'h20;
frames[19][27][22] = 8'h00;
frames[19][27][23] = 8'h00;
frames[19][27][24] = 8'h00;
frames[19][27][25] = 8'h00;
frames[19][27][26] = 8'h48;
frames[19][27][27] = 8'h6d;
frames[19][27][28] = 8'h92;
frames[19][27][29] = 8'h92;
frames[19][27][30] = 8'h92;
frames[19][27][31] = 8'h92;
frames[19][27][32] = 8'h92;
frames[19][27][33] = 8'h49;
frames[19][27][34] = 8'h6d;
frames[19][27][35] = 8'h92;
frames[19][27][36] = 8'h92;
frames[19][27][37] = 8'h6d;
frames[19][27][38] = 8'h24;
frames[19][27][39] = 8'h00;
frames[19][28][0] = 8'h24;
frames[19][28][1] = 8'h24;
frames[19][28][2] = 8'h24;
frames[19][28][3] = 8'h24;
frames[19][28][4] = 8'h24;
frames[19][28][5] = 8'h24;
frames[19][28][6] = 8'h24;
frames[19][28][7] = 8'h24;
frames[19][28][8] = 8'h24;
frames[19][28][9] = 8'h24;
frames[19][28][10] = 8'h24;
frames[19][28][11] = 8'h24;
frames[19][28][12] = 8'h24;
frames[19][28][13] = 8'h24;
frames[19][28][14] = 8'h24;
frames[19][28][15] = 8'h24;
frames[19][28][16] = 8'h24;
frames[19][28][17] = 8'h24;
frames[19][28][18] = 8'h20;
frames[19][28][19] = 8'h00;
frames[19][28][20] = 8'h00;
frames[19][28][21] = 8'h20;
frames[19][28][22] = 8'h20;
frames[19][28][23] = 8'h00;
frames[19][28][24] = 8'h00;
frames[19][28][25] = 8'h20;
frames[19][28][26] = 8'h24;
frames[19][28][27] = 8'h49;
frames[19][28][28] = 8'h49;
frames[19][28][29] = 8'h49;
frames[19][28][30] = 8'h49;
frames[19][28][31] = 8'h49;
frames[19][28][32] = 8'h49;
frames[19][28][33] = 8'h24;
frames[19][28][34] = 8'h49;
frames[19][28][35] = 8'h49;
frames[19][28][36] = 8'h49;
frames[19][28][37] = 8'h69;
frames[19][28][38] = 8'h24;
frames[19][28][39] = 8'h00;
frames[19][29][0] = 8'h24;
frames[19][29][1] = 8'h24;
frames[19][29][2] = 8'h24;
frames[19][29][3] = 8'h20;
frames[19][29][4] = 8'h20;
frames[19][29][5] = 8'h20;
frames[19][29][6] = 8'h20;
frames[19][29][7] = 8'h20;
frames[19][29][8] = 8'h24;
frames[19][29][9] = 8'h24;
frames[19][29][10] = 8'h24;
frames[19][29][11] = 8'h24;
frames[19][29][12] = 8'h24;
frames[19][29][13] = 8'h24;
frames[19][29][14] = 8'h24;
frames[19][29][15] = 8'h24;
frames[19][29][16] = 8'h24;
frames[19][29][17] = 8'h24;
frames[19][29][18] = 8'h20;
frames[19][29][19] = 8'h00;
frames[19][29][20] = 8'h00;
frames[19][29][21] = 8'h00;
frames[19][29][22] = 8'h20;
frames[19][29][23] = 8'h20;
frames[19][29][24] = 8'h00;
frames[19][29][25] = 8'h24;
frames[19][29][26] = 8'h24;
frames[19][29][27] = 8'h24;
frames[19][29][28] = 8'h00;
frames[19][29][29] = 8'h00;
frames[19][29][30] = 8'h00;
frames[19][29][31] = 8'h00;
frames[19][29][32] = 8'h00;
frames[19][29][33] = 8'h00;
frames[19][29][34] = 8'h00;
frames[19][29][35] = 8'h00;
frames[19][29][36] = 8'h00;
frames[19][29][37] = 8'h00;
frames[19][29][38] = 8'h24;
frames[19][29][39] = 8'h00;
	end
endmodule
